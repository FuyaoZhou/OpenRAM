VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_16x2
   CLASS BLOCK ;
   SIZE 464.48 BY 446.65 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  82.28 0.0 82.66 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  88.12 0.0 88.5 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.96 0.0 94.34 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.8 0.0 100.18 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.64 0.0 106.02 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  111.48 0.0 111.86 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  117.32 0.0 117.7 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.16 0.0 123.54 0.38 ;
      END
   END din0[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  64.76 0.0 65.14 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.6 0.0 70.98 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  76.44 0.0 76.82 0.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.185 0.38 143.565 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 151.585 0.38 151.965 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.79 0.38 158.17 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 166.29 0.38 166.67 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 171.93 0.38 172.31 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 180.43 0.38 180.81 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 186.675 0.38 187.055 ;
      END
   END addr0[9]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  394.88 446.27 395.26 446.65 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  389.04 446.27 389.42 446.65 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  383.2 446.27 383.58 446.65 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 98.51 464.48 98.89 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 90.01 464.48 90.39 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 84.37 464.48 84.75 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 75.87 464.48 76.25 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 70.23 464.48 70.61 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 61.73 464.48 62.11 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 56.09 464.48 56.47 ;
      END
   END addr1[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 42.385 0.38 42.765 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 398.3 464.48 398.68 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 50.785 0.38 51.165 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 43.875 0.38 44.255 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  464.1 397.555 464.48 397.935 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  133.265 0.0 133.645 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  158.225 0.0 158.605 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  183.185 0.0 183.565 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.145 0.0 208.525 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.105 0.0 233.485 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  258.065 0.0 258.445 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  283.025 0.0 283.405 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.985 0.0 308.365 0.38 ;
      END
   END dout0[7]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  133.325 446.27 133.705 446.65 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  158.285 446.27 158.665 446.65 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  183.245 446.27 183.625 446.65 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.205 446.27 208.585 446.65 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.165 446.27 233.545 446.65 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  258.125 446.27 258.505 446.65 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  283.085 446.27 283.465 446.65 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  308.045 446.27 308.425 446.65 ;
      END
   END dout1[7]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 446.65 ;
         LAYER met4 ;
         RECT  462.74 0.0 464.48 446.65 ;
         LAYER met3 ;
         RECT  0.0 444.91 464.48 446.65 ;
         LAYER met3 ;
         RECT  0.0 0.0 464.48 1.74 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.48 441.43 461.0 443.17 ;
         LAYER met4 ;
         RECT  459.26 3.48 461.0 443.17 ;
         LAYER met3 ;
         RECT  3.48 3.48 461.0 5.22 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 443.17 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 463.86 446.03 ;
   LAYER  met2 ;
      RECT  0.62 0.62 463.86 446.03 ;
   LAYER  met3 ;
      RECT  0.98 142.585 463.86 144.165 ;
      RECT  0.62 144.165 0.98 150.985 ;
      RECT  0.62 152.565 0.98 157.19 ;
      RECT  0.62 158.77 0.98 165.69 ;
      RECT  0.62 167.27 0.98 171.33 ;
      RECT  0.62 172.91 0.98 179.83 ;
      RECT  0.62 181.41 0.98 186.075 ;
      RECT  0.98 97.91 463.5 99.49 ;
      RECT  0.98 99.49 463.5 142.585 ;
      RECT  463.5 99.49 463.86 142.585 ;
      RECT  463.5 90.99 463.86 97.91 ;
      RECT  463.5 85.35 463.86 89.41 ;
      RECT  463.5 76.85 463.86 83.77 ;
      RECT  463.5 71.21 463.86 75.27 ;
      RECT  463.5 62.71 463.86 69.63 ;
      RECT  463.5 57.07 463.86 61.13 ;
      RECT  0.98 144.165 463.5 397.7 ;
      RECT  0.98 397.7 463.5 399.28 ;
      RECT  0.62 51.765 0.98 142.585 ;
      RECT  0.62 44.855 0.98 50.185 ;
      RECT  463.5 144.165 463.86 396.955 ;
      RECT  0.62 187.655 0.98 444.31 ;
      RECT  463.5 399.28 463.86 444.31 ;
      RECT  463.5 2.34 463.86 55.49 ;
      RECT  0.62 2.34 0.98 41.785 ;
      RECT  0.98 399.28 2.88 440.83 ;
      RECT  0.98 440.83 2.88 443.77 ;
      RECT  0.98 443.77 2.88 444.31 ;
      RECT  2.88 399.28 461.6 440.83 ;
      RECT  2.88 443.77 461.6 444.31 ;
      RECT  461.6 399.28 463.5 440.83 ;
      RECT  461.6 440.83 463.5 443.77 ;
      RECT  461.6 443.77 463.5 444.31 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 97.91 ;
      RECT  2.88 2.34 461.6 2.88 ;
      RECT  2.88 5.82 461.6 97.91 ;
      RECT  461.6 2.34 463.5 2.88 ;
      RECT  461.6 2.88 463.5 5.82 ;
      RECT  461.6 5.82 463.5 97.91 ;
   LAYER  met4 ;
      RECT  81.68 0.98 83.26 446.03 ;
      RECT  83.26 0.62 87.52 0.98 ;
      RECT  89.1 0.62 93.36 0.98 ;
      RECT  94.94 0.62 99.2 0.98 ;
      RECT  100.78 0.62 105.04 0.98 ;
      RECT  106.62 0.62 110.88 0.98 ;
      RECT  112.46 0.62 116.72 0.98 ;
      RECT  118.3 0.62 122.56 0.98 ;
      RECT  65.74 0.62 70.0 0.98 ;
      RECT  71.58 0.62 75.84 0.98 ;
      RECT  77.42 0.62 81.68 0.98 ;
      RECT  83.26 0.98 394.28 445.67 ;
      RECT  394.28 0.98 395.86 445.67 ;
      RECT  390.02 445.67 394.28 446.03 ;
      RECT  384.18 445.67 388.44 446.03 ;
      RECT  124.14 0.62 132.665 0.98 ;
      RECT  134.245 0.62 157.625 0.98 ;
      RECT  159.205 0.62 182.585 0.98 ;
      RECT  184.165 0.62 207.545 0.98 ;
      RECT  209.125 0.62 232.505 0.98 ;
      RECT  234.085 0.62 257.465 0.98 ;
      RECT  259.045 0.62 282.425 0.98 ;
      RECT  284.005 0.62 307.385 0.98 ;
      RECT  83.26 445.67 132.725 446.03 ;
      RECT  134.305 445.67 157.685 446.03 ;
      RECT  159.265 445.67 182.645 446.03 ;
      RECT  184.225 445.67 207.605 446.03 ;
      RECT  209.185 445.67 232.565 446.03 ;
      RECT  234.145 445.67 257.525 446.03 ;
      RECT  259.105 445.67 282.485 446.03 ;
      RECT  284.065 445.67 307.445 446.03 ;
      RECT  309.025 445.67 382.6 446.03 ;
      RECT  2.34 0.62 64.16 0.98 ;
      RECT  395.86 445.67 462.14 446.03 ;
      RECT  308.965 0.62 462.14 0.98 ;
      RECT  395.86 0.98 458.66 2.88 ;
      RECT  395.86 2.88 458.66 443.77 ;
      RECT  395.86 443.77 458.66 445.67 ;
      RECT  458.66 0.98 461.6 2.88 ;
      RECT  458.66 443.77 461.6 445.67 ;
      RECT  461.6 0.98 462.14 2.88 ;
      RECT  461.6 2.88 462.14 443.77 ;
      RECT  461.6 443.77 462.14 445.67 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 443.77 ;
      RECT  2.34 443.77 2.88 446.03 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 443.77 5.82 446.03 ;
      RECT  5.82 0.98 81.68 2.88 ;
      RECT  5.82 2.88 81.68 443.77 ;
      RECT  5.82 443.77 81.68 446.03 ;
   END
END    sky130_16x2
END    LIBRARY
