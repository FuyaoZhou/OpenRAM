**************************************************
* OpenRAM generated memory.
* Words: 256
* Data bits: 8
* Banks: 1
* Column mux: 8:1
* Trimmed: True
* LVS: False
**************************************************

* spice ptx M{0} {1} n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

* spice ptx M{0} {1} p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

* spice ptx M{0} {1} n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

* spice ptx M{0} {1} n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

.SUBCKT scn4m_subm_256x8_pnand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand3_pmos1 vdd A Z vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pnand3_0

* spice ptx M{0} {1} p m=2 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p

* spice ptx M{0} {1} n m=2 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p

.SUBCKT scn4m_subm_256x8_pinv_13
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 8
Mpinv_pmos Z A vdd vdd p m=2 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
Mpinv_nmos Z A gnd gnd n m=2 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
.ENDS scn4m_subm_256x8_pinv_13

.SUBCKT scn4m_subm_256x8_pdriver_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [8]
Xbuf_inv1
+ A Z vdd gnd
+ scn4m_subm_256x8_pinv_13
.ENDS scn4m_subm_256x8_pdriver_4

.SUBCKT scn4m_subm_256x8_pand3_1
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 8
Xpand3_nand
+ A B C zb_int vdd gnd
+ scn4m_subm_256x8_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pdriver_4
.ENDS scn4m_subm_256x8_pand3_1

* spice ptx M{0} {1} n m=4 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p

* spice ptx M{0} {1} p m=4 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p

.SUBCKT scn4m_subm_256x8_pinv_12
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 16
Mpinv_pmos Z A vdd vdd p m=4 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
Mpinv_nmos Z A gnd gnd n m=4 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
.ENDS scn4m_subm_256x8_pinv_12

.SUBCKT scn4m_subm_256x8_pdriver_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [16]
Xbuf_inv1
+ A Z vdd gnd
+ scn4m_subm_256x8_pinv_12
.ENDS scn4m_subm_256x8_pdriver_3

.SUBCKT scn4m_subm_256x8_pand3_0
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 16
Xpand3_nand
+ A B C zb_int vdd gnd
+ scn4m_subm_256x8_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pdriver_3
.ENDS scn4m_subm_256x8_pand3_0

* spice ptx M{0} {1} p m=5 w=6.7u l=0.4u pd=14.20u ps=14.20u as=6.70p ad=6.70p

* spice ptx M{0} {1} n m=5 w=3.4000000000000004u l=0.4u pd=7.60u ps=7.60u as=3.40p ad=3.40p

.SUBCKT scn4m_subm_256x8_pinv_16
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 21
Mpinv_pmos Z A vdd vdd p m=5 w=6.7u l=0.4u pd=14.20u ps=14.20u as=6.70p ad=6.70p
Mpinv_nmos Z A gnd gnd n m=5 w=3.4000000000000004u l=0.4u pd=7.60u ps=7.60u as=3.40p ad=3.40p
.ENDS scn4m_subm_256x8_pinv_16

* spice ptx M{0} {1} p m=1 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p

* spice ptx M{0} {1} n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

.SUBCKT scn4m_subm_256x8_pinv_14
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 2
Mpinv_pmos Z A vdd vdd p m=1 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
Mpinv_nmos Z A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pinv_14

* spice ptx M{0} {1} n m=2 w=2.8000000000000003u l=0.4u pd=6.40u ps=6.40u as=2.80p ad=2.80p

* spice ptx M{0} {1} p m=2 w=5.6000000000000005u l=0.4u pd=12.00u ps=12.00u as=5.60p ad=5.60p

.SUBCKT scn4m_subm_256x8_pinv_15
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 7
Mpinv_pmos Z A vdd vdd p m=2 w=5.6000000000000005u l=0.4u pd=12.00u ps=12.00u as=5.60p ad=5.60p
Mpinv_nmos Z A gnd gnd n m=2 w=2.8000000000000003u l=0.4u pd=6.40u ps=6.40u as=2.80p ad=2.80p
.ENDS scn4m_subm_256x8_pinv_15

* spice ptx M{0} {1} p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

* spice ptx M{0} {1} n m=1 w=0.8u l=0.4u pd=2.40u ps=2.40u as=0.80p ad=0.80p

.SUBCKT scn4m_subm_256x8_pinv_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpinv_nmos Z A gnd gnd n m=1 w=0.8u l=0.4u pd=2.40u ps=2.40u as=0.80p ad=0.80p
.ENDS scn4m_subm_256x8_pinv_1

.SUBCKT scn4m_subm_256x8_pdriver_5
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 2, 7, 21]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ scn4m_subm_256x8_pinv_1
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ scn4m_subm_256x8_pinv_14
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ scn4m_subm_256x8_pinv_15
Xbuf_inv4
+ Zb3_int Z vdd gnd
+ scn4m_subm_256x8_pinv_16
.ENDS scn4m_subm_256x8_pdriver_5

.SUBCKT scn4m_subm_256x8_pnand2_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand2_pmos1 vdd A Z vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pnand2_0

* spice ptx M{0} {1} n m=3 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p

* spice ptx M{0} {1} p m=3 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p

.SUBCKT scn4m_subm_256x8_pinv_5
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 12
Mpinv_pmos Z A vdd vdd p m=3 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
Mpinv_nmos Z A gnd gnd n m=3 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
.ENDS scn4m_subm_256x8_pinv_5

.SUBCKT scn4m_subm_256x8_pdriver_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [12]
Xbuf_inv1
+ A Z vdd gnd
+ scn4m_subm_256x8_pinv_5
.ENDS scn4m_subm_256x8_pdriver_0

.SUBCKT scn4m_subm_256x8_pand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 12
Xpand2_nand
+ A B zb_int vdd gnd
+ scn4m_subm_256x8_pnand2_0
Xpand2_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pdriver_0
.ENDS scn4m_subm_256x8_pand2

* spice ptx M{0} {1} p m=8 w=7.4u l=0.4u pd=15.60u ps=15.60u as=7.40p ad=7.40p

* spice ptx M{0} {1} n m=8 w=3.7u l=0.4u pd=8.20u ps=8.20u as=3.70p ad=3.70p

.SUBCKT scn4m_subm_256x8_pinv_9
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 37
Mpinv_pmos Z A vdd vdd p m=8 w=7.4u l=0.4u pd=15.60u ps=15.60u as=7.40p ad=7.40p
Mpinv_nmos Z A gnd gnd n m=8 w=3.7u l=0.4u pd=8.20u ps=8.20u as=3.70p ad=3.70p
.ENDS scn4m_subm_256x8_pinv_9

* spice ptx M{0} {1} p m=1 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p

* spice ptx M{0} {1} n m=1 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p

.SUBCKT scn4m_subm_256x8_pinv_8
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 4
Mpinv_pmos Z A vdd vdd p m=1 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
Mpinv_nmos Z A gnd gnd n m=1 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
.ENDS scn4m_subm_256x8_pinv_8

.SUBCKT scn4m_subm_256x8_pdriver_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 4, 12, 37]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ scn4m_subm_256x8_pinv_1
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ scn4m_subm_256x8_pinv_1
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ scn4m_subm_256x8_pinv_1
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ scn4m_subm_256x8_pinv_8
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ scn4m_subm_256x8_pinv_5
Xbuf_inv6
+ Zb5_int Z vdd gnd
+ scn4m_subm_256x8_pinv_9
.ENDS scn4m_subm_256x8_pdriver_1

.SUBCKT scn4m_subm_256x8_pinv_17
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpinv_nmos Z A gnd gnd n m=1 w=0.8u l=0.4u pd=2.40u ps=2.40u as=0.80p ad=0.80p
.ENDS scn4m_subm_256x8_pinv_17

.SUBCKT scn4m_subm_256x8_delay_chain
+ in out vdd gnd
* INPUT : in 
* OUTPUT: out 
* POWER : vdd 
* GROUND: gnd 
* fanouts: [4, 4, 4, 4, 4, 4, 4, 4, 4]
Xdinv0
+ in dout_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_0_0
+ dout_1 n_0_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_0_1
+ dout_1 n_0_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_0_2
+ dout_1 n_0_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_0_3
+ dout_1 n_0_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv1
+ dout_1 dout_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_1_0
+ dout_2 n_1_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_1_1
+ dout_2 n_1_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_1_2
+ dout_2 n_1_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_1_3
+ dout_2 n_1_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv2
+ dout_2 dout_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_2_0
+ dout_3 n_2_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_2_1
+ dout_3 n_2_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_2_2
+ dout_3 n_2_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_2_3
+ dout_3 n_2_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv3
+ dout_3 dout_4 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_3_0
+ dout_4 n_3_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_3_1
+ dout_4 n_3_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_3_2
+ dout_4 n_3_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_3_3
+ dout_4 n_3_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv4
+ dout_4 dout_5 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_4_0
+ dout_5 n_4_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_4_1
+ dout_5 n_4_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_4_2
+ dout_5 n_4_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_4_3
+ dout_5 n_4_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv5
+ dout_5 dout_6 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_5_0
+ dout_6 n_5_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_5_1
+ dout_6 n_5_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_5_2
+ dout_6 n_5_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_5_3
+ dout_6 n_5_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv6
+ dout_6 dout_7 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_6_0
+ dout_7 n_6_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_6_1
+ dout_7 n_6_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_6_2
+ dout_7 n_6_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_6_3
+ dout_7 n_6_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv7
+ dout_7 dout_8 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_7_0
+ dout_8 n_7_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_7_1
+ dout_8 n_7_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_7_2
+ dout_8 n_7_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_7_3
+ dout_8 n_7_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdinv8
+ dout_8 out vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_8_0
+ out n_8_0 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_8_1
+ out n_8_1 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_8_2
+ out n_8_2 vdd gnd
+ scn4m_subm_256x8_pinv_17
Xdload_8_3
+ out n_8_3 vdd gnd
+ scn4m_subm_256x8_pinv_17
.ENDS scn4m_subm_256x8_delay_chain

.SUBCKT scn4m_subm_256x8_pinv_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 4
Mpinv_pmos Z A vdd vdd p m=1 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
Mpinv_nmos Z A gnd gnd n m=1 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
.ENDS scn4m_subm_256x8_pinv_4
*********************** "dff" ******************************
* Positive edge-triggered FF
.SUBCKT dff D Q clk vdd gnd

* SPICE3 file created from dff.ext - technology: scmos

M1000 vdd clk a_24_24# vdd p w=8u l=0.4u
M1001 a_84_296# D vdd vdd p w=4u l=0.4u
M1002 a_104_24# clk a_84_296# vdd p w=4u l=0.4u
M1003 a_140_296# a_24_24# a_104_24# vdd p w=4u l=0.4u
M1004 vdd a_152_16# a_140_296# vdd p w=4u l=0.4u
M1005 a_152_16# a_104_24# vdd vdd p w=4u l=0.4u
M1006 a_260_296# a_152_16# vdd vdd p w=4u l=0.4u
M1007 a_280_24# a_24_24# a_260_296# vdd p w=4u l=0.4u
M1008 a_320_336# clk a_280_24# vdd p w=2u l=0.4u
M1009 vdd Q a_320_336# vdd p w=2u l=0.4u
M1010 gnd clk a_24_24# gnd n w=4u l=0.4u
M1011 Q a_280_24# vdd vdd p w=8u l=0.4u
M1012 a_84_24# D gnd gnd n w=2u l=0.4u
M1013 a_104_24# a_24_24# a_84_24# gnd n w=2u l=0.4u
M1014 a_140_24# clk a_104_24# gnd n w=2u l=0.4u
M1015 gnd a_152_16# a_140_24# gnd n w=2u l=0.4u
M1016 a_152_16# a_104_24# gnd gnd n w=2u l=0.4u
M1017 a_260_24# a_152_16# gnd gnd n w=2u l=0.4u
M1018 a_280_24# clk a_260_24# gnd n w=2u l=0.4u
M1019 a_320_24# a_24_24# a_280_24# gnd n w=2u l=0.4u
M1020 gnd Q a_320_24# gnd n w=2u l=0.4u
M1021 Q a_280_24# gnd gnd n w=4u l=0.4u

.ENDS

.SUBCKT scn4m_subm_256x8_pinv_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 2
Mpinv_pmos Z A vdd vdd p m=1 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
Mpinv_nmos Z A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pinv_3

.SUBCKT scn4m_subm_256x8_dff_buf_0
+ D Q Qb clk vdd gnd
* INPUT : D 
* OUTPUT: Q 
* OUTPUT: Qb 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* inv1: 2 inv2: 4
Xdff_buf_dff
+ D qint clk vdd gnd
+ dff
Xdff_buf_inv1
+ qint Qb vdd gnd
+ scn4m_subm_256x8_pinv_3
Xdff_buf_inv2
+ Qb Q vdd gnd
+ scn4m_subm_256x8_pinv_4
.ENDS scn4m_subm_256x8_dff_buf_0

.SUBCKT scn4m_subm_256x8_dff_buf_array
+ din_0 din_1 dout_0 dout_bar_0 dout_1 dout_bar_1 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* OUTPUT: dout_0 
* OUTPUT: dout_bar_0 
* OUTPUT: dout_1 
* OUTPUT: dout_bar_1 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 2 cols: 1
* inv1: 2 inv2: 4
Xdff_r0_c0
+ din_0 dout_0 dout_bar_0 clk vdd gnd
+ scn4m_subm_256x8_dff_buf_0
Xdff_r1_c0
+ din_1 dout_1 dout_bar_1 clk vdd gnd
+ scn4m_subm_256x8_dff_buf_0
.ENDS scn4m_subm_256x8_dff_buf_array

.SUBCKT scn4m_subm_256x8_pnand2_1
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand2_pmos1 vdd A Z vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pnand2_1

* spice ptx M{0} {1} p m=2 w=8.0u l=0.4u pd=16.80u ps=16.80u as=8.00p ad=8.00p

* spice ptx M{0} {1} n m=2 w=4.0u l=0.4u pd=8.80u ps=8.80u as=4.00p ad=4.00p

.SUBCKT scn4m_subm_256x8_pinv_11
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 10
Mpinv_pmos Z A vdd vdd p m=2 w=8.0u l=0.4u pd=16.80u ps=16.80u as=8.00p ad=8.00p
Mpinv_nmos Z A gnd gnd n m=2 w=4.0u l=0.4u pd=8.80u ps=8.80u as=4.00p ad=4.00p
.ENDS scn4m_subm_256x8_pinv_11

* spice ptx M{0} {1} n m=1 w=2.4000000000000004u l=0.4u pd=5.60u ps=5.60u as=2.40p ad=2.40p

* spice ptx M{0} {1} p m=1 w=4.800000000000001u l=0.4u pd=10.40u ps=10.40u as=4.80p ad=4.80p

.SUBCKT scn4m_subm_256x8_pinv_10
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 3
Mpinv_pmos Z A vdd vdd p m=1 w=4.800000000000001u l=0.4u pd=10.40u ps=10.40u as=4.80p ad=4.80p
Mpinv_nmos Z A gnd gnd n m=1 w=2.4000000000000004u l=0.4u pd=5.60u ps=5.60u as=2.40p ad=2.40p
.ENDS scn4m_subm_256x8_pinv_10

.SUBCKT scn4m_subm_256x8_pdriver_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [3, 10]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ scn4m_subm_256x8_pinv_10
Xbuf_inv2
+ Zb1_int Z vdd gnd
+ scn4m_subm_256x8_pinv_11
.ENDS scn4m_subm_256x8_pdriver_2

.SUBCKT scn4m_subm_256x8_pinv_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpinv_nmos Z A gnd gnd n m=1 w=0.8u l=0.4u pd=2.40u ps=2.40u as=0.80p ad=0.80p
.ENDS scn4m_subm_256x8_pinv_2

.SUBCKT scn4m_subm_256x8_control_logic_rw
+ csb web clk rbl_bl s_en w_en p_en_bar wl_en clk_buf vdd gnd
* INPUT : csb 
* INPUT : web 
* INPUT : clk 
* INPUT : rbl_bl 
* OUTPUT: s_en 
* OUTPUT: w_en 
* OUTPUT: p_en_bar 
* OUTPUT: wl_en 
* OUTPUT: clk_buf 
* POWER : vdd 
* GROUND: gnd 
* num_rows: 32
* words_per_row: 8
* word_size 8
Xctrl_dffs
+ csb web cs_bar cs we_bar we clk_buf vdd gnd
+ scn4m_subm_256x8_dff_buf_array
Xclkbuf
+ clk clk_buf vdd gnd
+ scn4m_subm_256x8_pdriver_1
Xinv_clk_bar
+ clk_buf clk_bar vdd gnd
+ scn4m_subm_256x8_pinv_2
Xand2_gated_clk_bar
+ clk_bar cs gated_clk_bar vdd gnd
+ scn4m_subm_256x8_pand2
Xand2_gated_clk_buf
+ clk_buf cs gated_clk_buf vdd gnd
+ scn4m_subm_256x8_pand2
Xbuf_wl_en
+ gated_clk_bar wl_en vdd gnd
+ scn4m_subm_256x8_pdriver_2
Xrbl_bl_delay_inv
+ rbl_bl_delay rbl_bl_delay_bar vdd gnd
+ scn4m_subm_256x8_pinv_2
Xw_en_and
+ we rbl_bl_delay_bar gated_clk_bar w_en vdd gnd
+ scn4m_subm_256x8_pand3_0
Xbuf_s_en_and
+ rbl_bl_delay gated_clk_bar we_bar s_en vdd gnd
+ scn4m_subm_256x8_pand3_1
Xdelay_chain
+ rbl_bl rbl_bl_delay vdd gnd
+ scn4m_subm_256x8_delay_chain
Xnand_p_en_bar
+ gated_clk_buf rbl_bl_delay p_en_bar_unbuf vdd gnd
+ scn4m_subm_256x8_pnand2_1
Xbuf_p_en_bar
+ p_en_bar_unbuf p_en_bar vdd gnd
+ scn4m_subm_256x8_pdriver_5
.ENDS scn4m_subm_256x8_control_logic_rw

* spice ptx M{0} {1} n m=1 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p

.SUBCKT scn4m_subm_256x8_column_mux
+ bl br bl_out br_out sel gnd
* INOUT : bl 
* INOUT : br 
* INOUT : bl_out 
* INOUT : br_out 
* INOUT : sel 
* INOUT : gnd 
Mmux_tx1 bl sel bl_out gnd n m=1 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
Mmux_tx2 br sel br_out gnd n m=1 w=6.4u l=0.4u pd=13.60u ps=13.60u as=6.40p ad=6.40p
.ENDS scn4m_subm_256x8_column_mux

.SUBCKT scn4m_subm_256x8_column_mux_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7
+ bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3
+ br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6
+ bl_out_7 br_out_7 gnd
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : sel_2 
* INOUT : sel_3 
* INOUT : sel_4 
* INOUT : sel_5 
* INOUT : sel_6 
* INOUT : sel_7 
* INOUT : bl_out_0 
* INOUT : br_out_0 
* INOUT : bl_out_1 
* INOUT : br_out_1 
* INOUT : bl_out_2 
* INOUT : br_out_2 
* INOUT : bl_out_3 
* INOUT : br_out_3 
* INOUT : bl_out_4 
* INOUT : br_out_4 
* INOUT : bl_out_5 
* INOUT : br_out_5 
* INOUT : bl_out_6 
* INOUT : br_out_6 
* INOUT : bl_out_7 
* INOUT : br_out_7 
* INOUT : gnd 
* cols: 64 word_size: 8 bl: bl br: br
XXMUX0
+ bl_0 br_0 bl_out_0 br_out_0 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX1
+ bl_1 br_1 bl_out_0 br_out_0 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX2
+ bl_2 br_2 bl_out_0 br_out_0 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX3
+ bl_3 br_3 bl_out_0 br_out_0 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX4
+ bl_4 br_4 bl_out_0 br_out_0 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX5
+ bl_5 br_5 bl_out_0 br_out_0 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX6
+ bl_6 br_6 bl_out_0 br_out_0 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX7
+ bl_7 br_7 bl_out_0 br_out_0 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX8
+ bl_8 br_8 bl_out_1 br_out_1 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX9
+ bl_9 br_9 bl_out_1 br_out_1 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX10
+ bl_10 br_10 bl_out_1 br_out_1 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX11
+ bl_11 br_11 bl_out_1 br_out_1 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX12
+ bl_12 br_12 bl_out_1 br_out_1 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX13
+ bl_13 br_13 bl_out_1 br_out_1 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX14
+ bl_14 br_14 bl_out_1 br_out_1 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX15
+ bl_15 br_15 bl_out_1 br_out_1 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX16
+ bl_16 br_16 bl_out_2 br_out_2 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX17
+ bl_17 br_17 bl_out_2 br_out_2 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX18
+ bl_18 br_18 bl_out_2 br_out_2 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX19
+ bl_19 br_19 bl_out_2 br_out_2 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX20
+ bl_20 br_20 bl_out_2 br_out_2 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX21
+ bl_21 br_21 bl_out_2 br_out_2 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX22
+ bl_22 br_22 bl_out_2 br_out_2 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX23
+ bl_23 br_23 bl_out_2 br_out_2 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX24
+ bl_24 br_24 bl_out_3 br_out_3 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX25
+ bl_25 br_25 bl_out_3 br_out_3 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX26
+ bl_26 br_26 bl_out_3 br_out_3 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX27
+ bl_27 br_27 bl_out_3 br_out_3 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX28
+ bl_28 br_28 bl_out_3 br_out_3 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX29
+ bl_29 br_29 bl_out_3 br_out_3 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX30
+ bl_30 br_30 bl_out_3 br_out_3 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX31
+ bl_31 br_31 bl_out_3 br_out_3 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX32
+ bl_32 br_32 bl_out_4 br_out_4 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX33
+ bl_33 br_33 bl_out_4 br_out_4 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX34
+ bl_34 br_34 bl_out_4 br_out_4 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX35
+ bl_35 br_35 bl_out_4 br_out_4 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX36
+ bl_36 br_36 bl_out_4 br_out_4 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX37
+ bl_37 br_37 bl_out_4 br_out_4 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX38
+ bl_38 br_38 bl_out_4 br_out_4 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX39
+ bl_39 br_39 bl_out_4 br_out_4 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX40
+ bl_40 br_40 bl_out_5 br_out_5 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX41
+ bl_41 br_41 bl_out_5 br_out_5 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX42
+ bl_42 br_42 bl_out_5 br_out_5 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX43
+ bl_43 br_43 bl_out_5 br_out_5 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX44
+ bl_44 br_44 bl_out_5 br_out_5 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX45
+ bl_45 br_45 bl_out_5 br_out_5 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX46
+ bl_46 br_46 bl_out_5 br_out_5 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX47
+ bl_47 br_47 bl_out_5 br_out_5 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX48
+ bl_48 br_48 bl_out_6 br_out_6 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX49
+ bl_49 br_49 bl_out_6 br_out_6 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX50
+ bl_50 br_50 bl_out_6 br_out_6 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX51
+ bl_51 br_51 bl_out_6 br_out_6 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX52
+ bl_52 br_52 bl_out_6 br_out_6 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX53
+ bl_53 br_53 bl_out_6 br_out_6 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX54
+ bl_54 br_54 bl_out_6 br_out_6 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX55
+ bl_55 br_55 bl_out_6 br_out_6 sel_7 gnd
+ scn4m_subm_256x8_column_mux
XXMUX56
+ bl_56 br_56 bl_out_7 br_out_7 sel_0 gnd
+ scn4m_subm_256x8_column_mux
XXMUX57
+ bl_57 br_57 bl_out_7 br_out_7 sel_1 gnd
+ scn4m_subm_256x8_column_mux
XXMUX58
+ bl_58 br_58 bl_out_7 br_out_7 sel_2 gnd
+ scn4m_subm_256x8_column_mux
XXMUX59
+ bl_59 br_59 bl_out_7 br_out_7 sel_3 gnd
+ scn4m_subm_256x8_column_mux
XXMUX60
+ bl_60 br_60 bl_out_7 br_out_7 sel_4 gnd
+ scn4m_subm_256x8_column_mux
XXMUX61
+ bl_61 br_61 bl_out_7 br_out_7 sel_5 gnd
+ scn4m_subm_256x8_column_mux
XXMUX62
+ bl_62 br_62 bl_out_7 br_out_7 sel_6 gnd
+ scn4m_subm_256x8_column_mux
XXMUX63
+ bl_63 br_63 bl_out_7 br_out_7 sel_7 gnd
+ scn4m_subm_256x8_column_mux
.ENDS scn4m_subm_256x8_column_mux_array
*********************** "sense_amp" ******************************

.SUBCKT sense_amp bl br dout en vdd gnd

* SPICE3 file created from sense_amp.ext - technology: scmos

M1000 gnd en a_56_432# gnd n w=1.8u l=0.4u
M1001 a_56_432# a_48_304# dint gnd n w=1.8u l=0.4u
M1002 a_48_304# dint a_56_432# gnd n w=1.8u l=0.4u
M1003 vdd a_48_304# dint vdd p w=3.6u l=0.4u
M1004 a_48_304# dint vdd vdd p w=3.6u l=0.4u
M1005 bl en dint vdd p w=4.8u l=0.4u
M1006 a_48_304# en br vdd p w=4.8u l=0.4u

M1007 dout_bar dint vdd vdd p w=1.6u l=0.4u
M1008 gnd dint dout_bar gnd n w=0.8u l=0.4u
M1009 dout dout_bar vdd vdd p w=4.8u l=0.4u
M1010 gnd dout_bar dout gnd n w=2.4u l=0.4u
.ENDS

.SUBCKT scn4m_subm_256x8_sense_amp_array
+ data_0 bl_0 br_0 data_1 bl_1 br_1 data_2 bl_2 br_2 data_3 bl_3 br_3
+ data_4 bl_4 br_4 data_5 bl_5 br_5 data_6 bl_6 br_6 data_7 bl_7 br_7 en
+ vdd gnd
* OUTPUT: data_0 
* INPUT : bl_0 
* INPUT : br_0 
* OUTPUT: data_1 
* INPUT : bl_1 
* INPUT : br_1 
* OUTPUT: data_2 
* INPUT : bl_2 
* INPUT : br_2 
* OUTPUT: data_3 
* INPUT : bl_3 
* INPUT : br_3 
* OUTPUT: data_4 
* INPUT : bl_4 
* INPUT : br_4 
* OUTPUT: data_5 
* INPUT : bl_5 
* INPUT : br_5 
* OUTPUT: data_6 
* INPUT : bl_6 
* INPUT : br_6 
* OUTPUT: data_7 
* INPUT : bl_7 
* INPUT : br_7 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* word_size 8
* words_per_row: 8
Xsa_d0
+ bl_0 br_0 data_0 en vdd gnd
+ sense_amp
Xsa_d1
+ bl_1 br_1 data_1 en vdd gnd
+ sense_amp
Xsa_d2
+ bl_2 br_2 data_2 en vdd gnd
+ sense_amp
Xsa_d3
+ bl_3 br_3 data_3 en vdd gnd
+ sense_amp
Xsa_d4
+ bl_4 br_4 data_4 en vdd gnd
+ sense_amp
Xsa_d5
+ bl_5 br_5 data_5 en vdd gnd
+ sense_amp
Xsa_d6
+ bl_6 br_6 data_6 en vdd gnd
+ sense_amp
Xsa_d7
+ bl_7 br_7 data_7 en vdd gnd
+ sense_amp
.ENDS scn4m_subm_256x8_sense_amp_array
*********************** Write_Driver ******************************
.SUBCKT write_driver din bl br en vdd gnd

**** Inverter to conver Data_in to data_in_bar ******
* din_bar = inv(din)
M_1 din_bar din gnd gnd n W=0.8u L=0.4u
M_2 din_bar din vdd vdd p W=1.4u L=0.4u

**** 2input nand gate follwed by inverter to drive BL ******
* din_bar_gated = nand(en, din)
M_3 din_bar_gated en net_7 gnd n W=1.4u L=0.4u
M_4 net_7 din gnd gnd n W=1.4u L=0.4u
M_5 din_bar_gated en vdd vdd p W=1.4u L=0.4u
M_6 din_bar_gated din vdd vdd p W=1.4u L=0.4u
* din_bar_gated_bar = inv(din_bar_gated)
M_7 din_bar_gated_bar din_bar_gated vdd vdd p W=1.4u L=0.4u
M_8 din_bar_gated_bar din_bar_gated gnd gnd n W=0.8u L=0.4u

**** 2input nand gate follwed by inverter to drive BR******
* din_gated = nand(en, din_bar)
M_9 din_gated en vdd vdd p W=1.4u L=0.4u
M_10 din_gated en net_8 gnd n W=1.4u L=0.4u
M_11 net_8 din_bar gnd gnd n W=1.4u L=0.4u
M_12 din_gated din_bar vdd vdd p W=1.4u L=0.4u
* din_gated_bar = inv(din_gated)
M_13 din_gated_bar din_gated vdd vdd p W=1.4u L=0.4u
M_14 din_gated_bar din_gated gnd gnd n W=0.8u L=0.4u

************************************************
* pull down with en enable
M_15 bl din_gated_bar gnd gnd n W=2.4u L=0.4u
M_16 br din_bar_gated_bar gnd gnd n W=2.4u L=0.4u



.ENDS   $ write_driver

.SUBCKT scn4m_subm_256x8_write_driver_array
+ data_0 data_1 data_2 data_3 data_4 data_5 data_6 data_7 bl_0 br_0 bl_1
+ br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6 bl_7 br_7 en
+ vdd gnd
* INPUT : data_0 
* INPUT : data_1 
* INPUT : data_2 
* INPUT : data_3 
* INPUT : data_4 
* INPUT : data_5 
* INPUT : data_6 
* INPUT : data_7 
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* columns: 64
* word_size 8
Xwrite_driver0
+ data_0 bl_0 br_0 en vdd gnd
+ write_driver
Xwrite_driver8
+ data_1 bl_1 br_1 en vdd gnd
+ write_driver
Xwrite_driver16
+ data_2 bl_2 br_2 en vdd gnd
+ write_driver
Xwrite_driver24
+ data_3 bl_3 br_3 en vdd gnd
+ write_driver
Xwrite_driver32
+ data_4 bl_4 br_4 en vdd gnd
+ write_driver
Xwrite_driver40
+ data_5 bl_5 br_5 en vdd gnd
+ write_driver
Xwrite_driver48
+ data_6 bl_6 br_6 en vdd gnd
+ write_driver
Xwrite_driver56
+ data_7 bl_7 br_7 en vdd gnd
+ write_driver
.ENDS scn4m_subm_256x8_write_driver_array

.SUBCKT scn4m_subm_256x8_precharge_0
+ bl br en_bar vdd
* OUTPUT: bl 
* OUTPUT: br 
* INPUT : en_bar 
* POWER : vdd 
Mlower_pmos bl en_bar br vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mupper_pmos1 bl en_bar vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mupper_pmos2 br en_bar vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_precharge_0

.SUBCKT scn4m_subm_256x8_precharge_array
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 bl_64 br_64 en_bar vdd
* OUTPUT: bl_0 
* OUTPUT: br_0 
* OUTPUT: bl_1 
* OUTPUT: br_1 
* OUTPUT: bl_2 
* OUTPUT: br_2 
* OUTPUT: bl_3 
* OUTPUT: br_3 
* OUTPUT: bl_4 
* OUTPUT: br_4 
* OUTPUT: bl_5 
* OUTPUT: br_5 
* OUTPUT: bl_6 
* OUTPUT: br_6 
* OUTPUT: bl_7 
* OUTPUT: br_7 
* OUTPUT: bl_8 
* OUTPUT: br_8 
* OUTPUT: bl_9 
* OUTPUT: br_9 
* OUTPUT: bl_10 
* OUTPUT: br_10 
* OUTPUT: bl_11 
* OUTPUT: br_11 
* OUTPUT: bl_12 
* OUTPUT: br_12 
* OUTPUT: bl_13 
* OUTPUT: br_13 
* OUTPUT: bl_14 
* OUTPUT: br_14 
* OUTPUT: bl_15 
* OUTPUT: br_15 
* OUTPUT: bl_16 
* OUTPUT: br_16 
* OUTPUT: bl_17 
* OUTPUT: br_17 
* OUTPUT: bl_18 
* OUTPUT: br_18 
* OUTPUT: bl_19 
* OUTPUT: br_19 
* OUTPUT: bl_20 
* OUTPUT: br_20 
* OUTPUT: bl_21 
* OUTPUT: br_21 
* OUTPUT: bl_22 
* OUTPUT: br_22 
* OUTPUT: bl_23 
* OUTPUT: br_23 
* OUTPUT: bl_24 
* OUTPUT: br_24 
* OUTPUT: bl_25 
* OUTPUT: br_25 
* OUTPUT: bl_26 
* OUTPUT: br_26 
* OUTPUT: bl_27 
* OUTPUT: br_27 
* OUTPUT: bl_28 
* OUTPUT: br_28 
* OUTPUT: bl_29 
* OUTPUT: br_29 
* OUTPUT: bl_30 
* OUTPUT: br_30 
* OUTPUT: bl_31 
* OUTPUT: br_31 
* OUTPUT: bl_32 
* OUTPUT: br_32 
* OUTPUT: bl_33 
* OUTPUT: br_33 
* OUTPUT: bl_34 
* OUTPUT: br_34 
* OUTPUT: bl_35 
* OUTPUT: br_35 
* OUTPUT: bl_36 
* OUTPUT: br_36 
* OUTPUT: bl_37 
* OUTPUT: br_37 
* OUTPUT: bl_38 
* OUTPUT: br_38 
* OUTPUT: bl_39 
* OUTPUT: br_39 
* OUTPUT: bl_40 
* OUTPUT: br_40 
* OUTPUT: bl_41 
* OUTPUT: br_41 
* OUTPUT: bl_42 
* OUTPUT: br_42 
* OUTPUT: bl_43 
* OUTPUT: br_43 
* OUTPUT: bl_44 
* OUTPUT: br_44 
* OUTPUT: bl_45 
* OUTPUT: br_45 
* OUTPUT: bl_46 
* OUTPUT: br_46 
* OUTPUT: bl_47 
* OUTPUT: br_47 
* OUTPUT: bl_48 
* OUTPUT: br_48 
* OUTPUT: bl_49 
* OUTPUT: br_49 
* OUTPUT: bl_50 
* OUTPUT: br_50 
* OUTPUT: bl_51 
* OUTPUT: br_51 
* OUTPUT: bl_52 
* OUTPUT: br_52 
* OUTPUT: bl_53 
* OUTPUT: br_53 
* OUTPUT: bl_54 
* OUTPUT: br_54 
* OUTPUT: bl_55 
* OUTPUT: br_55 
* OUTPUT: bl_56 
* OUTPUT: br_56 
* OUTPUT: bl_57 
* OUTPUT: br_57 
* OUTPUT: bl_58 
* OUTPUT: br_58 
* OUTPUT: bl_59 
* OUTPUT: br_59 
* OUTPUT: bl_60 
* OUTPUT: br_60 
* OUTPUT: bl_61 
* OUTPUT: br_61 
* OUTPUT: bl_62 
* OUTPUT: br_62 
* OUTPUT: bl_63 
* OUTPUT: br_63 
* OUTPUT: bl_64 
* OUTPUT: br_64 
* INPUT : en_bar 
* POWER : vdd 
* cols: 65 size: 1 bl: bl br: br
Xpre_column_0
+ bl_0 br_0 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_1
+ bl_1 br_1 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_2
+ bl_2 br_2 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_3
+ bl_3 br_3 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_4
+ bl_4 br_4 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_5
+ bl_5 br_5 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_6
+ bl_6 br_6 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_7
+ bl_7 br_7 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_8
+ bl_8 br_8 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_9
+ bl_9 br_9 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_10
+ bl_10 br_10 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_11
+ bl_11 br_11 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_12
+ bl_12 br_12 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_13
+ bl_13 br_13 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_14
+ bl_14 br_14 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_15
+ bl_15 br_15 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_16
+ bl_16 br_16 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_17
+ bl_17 br_17 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_18
+ bl_18 br_18 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_19
+ bl_19 br_19 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_20
+ bl_20 br_20 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_21
+ bl_21 br_21 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_22
+ bl_22 br_22 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_23
+ bl_23 br_23 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_24
+ bl_24 br_24 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_25
+ bl_25 br_25 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_26
+ bl_26 br_26 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_27
+ bl_27 br_27 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_28
+ bl_28 br_28 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_29
+ bl_29 br_29 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_30
+ bl_30 br_30 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_31
+ bl_31 br_31 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_32
+ bl_32 br_32 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_33
+ bl_33 br_33 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_34
+ bl_34 br_34 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_35
+ bl_35 br_35 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_36
+ bl_36 br_36 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_37
+ bl_37 br_37 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_38
+ bl_38 br_38 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_39
+ bl_39 br_39 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_40
+ bl_40 br_40 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_41
+ bl_41 br_41 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_42
+ bl_42 br_42 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_43
+ bl_43 br_43 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_44
+ bl_44 br_44 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_45
+ bl_45 br_45 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_46
+ bl_46 br_46 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_47
+ bl_47 br_47 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_48
+ bl_48 br_48 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_49
+ bl_49 br_49 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_50
+ bl_50 br_50 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_51
+ bl_51 br_51 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_52
+ bl_52 br_52 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_53
+ bl_53 br_53 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_54
+ bl_54 br_54 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_55
+ bl_55 br_55 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_56
+ bl_56 br_56 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_57
+ bl_57 br_57 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_58
+ bl_58 br_58 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_59
+ bl_59 br_59 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_60
+ bl_60 br_60 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_61
+ bl_61 br_61 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_62
+ bl_62 br_62 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_63
+ bl_63 br_63 en_bar vdd
+ scn4m_subm_256x8_precharge_0
Xpre_column_64
+ bl_64 br_64 en_bar vdd
+ scn4m_subm_256x8_precharge_0
.ENDS scn4m_subm_256x8_precharge_array

.SUBCKT scn4m_subm_256x8_port_data
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 dout_0 dout_1 dout_2 dout_3 dout_4
+ dout_5 dout_6 dout_7 din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7
+ sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7 s_en p_en_bar w_en vdd
+ gnd
* INOUT : rbl_bl 
* INOUT : rbl_br 
* INOUT : bl_0 
* INOUT : br_0 
* INOUT : bl_1 
* INOUT : br_1 
* INOUT : bl_2 
* INOUT : br_2 
* INOUT : bl_3 
* INOUT : br_3 
* INOUT : bl_4 
* INOUT : br_4 
* INOUT : bl_5 
* INOUT : br_5 
* INOUT : bl_6 
* INOUT : br_6 
* INOUT : bl_7 
* INOUT : br_7 
* INOUT : bl_8 
* INOUT : br_8 
* INOUT : bl_9 
* INOUT : br_9 
* INOUT : bl_10 
* INOUT : br_10 
* INOUT : bl_11 
* INOUT : br_11 
* INOUT : bl_12 
* INOUT : br_12 
* INOUT : bl_13 
* INOUT : br_13 
* INOUT : bl_14 
* INOUT : br_14 
* INOUT : bl_15 
* INOUT : br_15 
* INOUT : bl_16 
* INOUT : br_16 
* INOUT : bl_17 
* INOUT : br_17 
* INOUT : bl_18 
* INOUT : br_18 
* INOUT : bl_19 
* INOUT : br_19 
* INOUT : bl_20 
* INOUT : br_20 
* INOUT : bl_21 
* INOUT : br_21 
* INOUT : bl_22 
* INOUT : br_22 
* INOUT : bl_23 
* INOUT : br_23 
* INOUT : bl_24 
* INOUT : br_24 
* INOUT : bl_25 
* INOUT : br_25 
* INOUT : bl_26 
* INOUT : br_26 
* INOUT : bl_27 
* INOUT : br_27 
* INOUT : bl_28 
* INOUT : br_28 
* INOUT : bl_29 
* INOUT : br_29 
* INOUT : bl_30 
* INOUT : br_30 
* INOUT : bl_31 
* INOUT : br_31 
* INOUT : bl_32 
* INOUT : br_32 
* INOUT : bl_33 
* INOUT : br_33 
* INOUT : bl_34 
* INOUT : br_34 
* INOUT : bl_35 
* INOUT : br_35 
* INOUT : bl_36 
* INOUT : br_36 
* INOUT : bl_37 
* INOUT : br_37 
* INOUT : bl_38 
* INOUT : br_38 
* INOUT : bl_39 
* INOUT : br_39 
* INOUT : bl_40 
* INOUT : br_40 
* INOUT : bl_41 
* INOUT : br_41 
* INOUT : bl_42 
* INOUT : br_42 
* INOUT : bl_43 
* INOUT : br_43 
* INOUT : bl_44 
* INOUT : br_44 
* INOUT : bl_45 
* INOUT : br_45 
* INOUT : bl_46 
* INOUT : br_46 
* INOUT : bl_47 
* INOUT : br_47 
* INOUT : bl_48 
* INOUT : br_48 
* INOUT : bl_49 
* INOUT : br_49 
* INOUT : bl_50 
* INOUT : br_50 
* INOUT : bl_51 
* INOUT : br_51 
* INOUT : bl_52 
* INOUT : br_52 
* INOUT : bl_53 
* INOUT : br_53 
* INOUT : bl_54 
* INOUT : br_54 
* INOUT : bl_55 
* INOUT : br_55 
* INOUT : bl_56 
* INOUT : br_56 
* INOUT : bl_57 
* INOUT : br_57 
* INOUT : bl_58 
* INOUT : br_58 
* INOUT : bl_59 
* INOUT : br_59 
* INOUT : bl_60 
* INOUT : br_60 
* INOUT : bl_61 
* INOUT : br_61 
* INOUT : bl_62 
* INOUT : br_62 
* INOUT : bl_63 
* INOUT : br_63 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* INPUT : sel_0 
* INPUT : sel_1 
* INPUT : sel_2 
* INPUT : sel_3 
* INPUT : sel_4 
* INPUT : sel_5 
* INPUT : sel_6 
* INPUT : sel_7 
* INPUT : s_en 
* INPUT : p_en_bar 
* INPUT : w_en 
* POWER : vdd 
* GROUND: gnd 
Xprecharge_array0
+ rbl_bl rbl_br bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5
+ br_5 bl_6 br_6 bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11
+ bl_12 br_12 bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17
+ br_17 bl_18 br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22
+ bl_23 br_23 bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28
+ br_28 bl_29 br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33
+ bl_34 br_34 bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39
+ br_39 bl_40 br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44
+ bl_45 br_45 bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50
+ br_50 bl_51 br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55
+ bl_56 br_56 bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61
+ br_61 bl_62 br_62 bl_63 br_63 p_en_bar vdd
+ scn4m_subm_256x8_precharge_array
Xsense_amp_array0
+ dout_0 bl_out_0 br_out_0 dout_1 bl_out_1 br_out_1 dout_2 bl_out_2
+ br_out_2 dout_3 bl_out_3 br_out_3 dout_4 bl_out_4 br_out_4 dout_5
+ bl_out_5 br_out_5 dout_6 bl_out_6 br_out_6 dout_7 bl_out_7 br_out_7
+ s_en vdd gnd
+ scn4m_subm_256x8_sense_amp_array
Xwrite_driver_array0
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 bl_out_0 br_out_0
+ bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3 br_out_3 bl_out_4
+ br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6 bl_out_7 br_out_7 w_en
+ vdd gnd
+ scn4m_subm_256x8_write_driver_array
Xcolumn_mux_array0
+ bl_0 br_0 bl_1 br_1 bl_2 br_2 bl_3 br_3 bl_4 br_4 bl_5 br_5 bl_6 br_6
+ bl_7 br_7 bl_8 br_8 bl_9 br_9 bl_10 br_10 bl_11 br_11 bl_12 br_12
+ bl_13 br_13 bl_14 br_14 bl_15 br_15 bl_16 br_16 bl_17 br_17 bl_18
+ br_18 bl_19 br_19 bl_20 br_20 bl_21 br_21 bl_22 br_22 bl_23 br_23
+ bl_24 br_24 bl_25 br_25 bl_26 br_26 bl_27 br_27 bl_28 br_28 bl_29
+ br_29 bl_30 br_30 bl_31 br_31 bl_32 br_32 bl_33 br_33 bl_34 br_34
+ bl_35 br_35 bl_36 br_36 bl_37 br_37 bl_38 br_38 bl_39 br_39 bl_40
+ br_40 bl_41 br_41 bl_42 br_42 bl_43 br_43 bl_44 br_44 bl_45 br_45
+ bl_46 br_46 bl_47 br_47 bl_48 br_48 bl_49 br_49 bl_50 br_50 bl_51
+ br_51 bl_52 br_52 bl_53 br_53 bl_54 br_54 bl_55 br_55 bl_56 br_56
+ bl_57 br_57 bl_58 br_58 bl_59 br_59 bl_60 br_60 bl_61 br_61 bl_62
+ br_62 bl_63 br_63 sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7
+ bl_out_0 br_out_0 bl_out_1 br_out_1 bl_out_2 br_out_2 bl_out_3
+ br_out_3 bl_out_4 br_out_4 bl_out_5 br_out_5 bl_out_6 br_out_6
+ bl_out_7 br_out_7 gnd
+ scn4m_subm_256x8_column_mux_array
.ENDS scn4m_subm_256x8_port_data

*********************** "dummy_cell_1rw" ******************************
.SUBCKT dummy_cell_1rw bl br wl vdd gnd

* Inverter 1
M1000 Q Q_bar vdd vdd p w=0.6u l=0.8u
M1002 Q Q_bar gnd gnd n w=1.6u l=0.4u

* Inverter 2
M1001 vdd Q Q_bar vdd p w=0.6u l=0.8u
M1003 gnd Q Q_bar gnd n w=1.6u l=0.4u

* Access transistors
M1004 Q wl bl_noconn gnd n w=0.8u l=0.4u
M1005 Q_bar wl br_noconn gnd n w=0.8u l=0.4u

.ENDS

.SUBCKT scn4m_subm_256x8_dummy_array_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS scn4m_subm_256x8_dummy_array_0

.SUBCKT scn4m_subm_256x8_dummy_array_2
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ dummy_cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ dummy_cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ dummy_cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ dummy_cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ dummy_cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ dummy_cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ dummy_cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ dummy_cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ dummy_cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ dummy_cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ dummy_cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ dummy_cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ dummy_cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ dummy_cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ dummy_cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ dummy_cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ dummy_cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ dummy_cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ dummy_cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ dummy_cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ dummy_cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ dummy_cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ dummy_cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ dummy_cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ dummy_cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ dummy_cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ dummy_cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ dummy_cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ dummy_cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ dummy_cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ dummy_cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ dummy_cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ dummy_cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ dummy_cell_1rw
.ENDS scn4m_subm_256x8_dummy_array_2

.SUBCKT scn4m_subm_256x8_dummy_array_3
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ dummy_cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ dummy_cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ dummy_cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ dummy_cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ dummy_cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ dummy_cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ dummy_cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ dummy_cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ dummy_cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ dummy_cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ dummy_cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ dummy_cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ dummy_cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ dummy_cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ dummy_cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ dummy_cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ dummy_cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ dummy_cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ dummy_cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ dummy_cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ dummy_cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ dummy_cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ dummy_cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ dummy_cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ dummy_cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ dummy_cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ dummy_cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ dummy_cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ dummy_cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ dummy_cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ dummy_cell_1rw
Xbit_r32_c0
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ dummy_cell_1rw
Xbit_r33_c0
+ bl_0_0 br_0_0 wl_0_33 vdd gnd
+ dummy_cell_1rw
Xbit_r34_c0
+ bl_0_0 br_0_0 wl_0_34 vdd gnd
+ dummy_cell_1rw
.ENDS scn4m_subm_256x8_dummy_array_3

.SUBCKT scn4m_subm_256x8_dummy_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS scn4m_subm_256x8_dummy_array

*********************** "cell_1rw" ******************************
.SUBCKT replica_cell_1rw bl br wl vdd gnd
* SPICE3 file created from cell_1rw.ext - technology: scmos

* Inverter 1
M1000 Q vdd vdd vdd p w=0.6u l=0.8u
M1002 Q vdd gnd gnd n w=1.6u l=0.4u

* Inverter 2
M1001 vdd Q vdd vdd p w=0.6u l=0.8u
M1003 gnd Q vdd gnd n w=1.6u l=0.4u

* Access transistors
M1004 Q wl bl gnd n w=0.8u l=0.4u
M1005 vdd wl br gnd n w=0.8u l=0.4u

.ENDS

.SUBCKT scn4m_subm_256x8_replica_column
+ bl_0_0 br_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32 vdd
+ gnd
* OUTPUT: bl_0_0 
* OUTPUT: br_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* POWER : vdd 
* GROUND: gnd 
Xrbc_0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ replica_cell_1rw
Xrbc_1
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ replica_cell_1rw
Xrbc_2
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ replica_cell_1rw
Xrbc_3
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ replica_cell_1rw
Xrbc_4
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ replica_cell_1rw
Xrbc_5
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ replica_cell_1rw
Xrbc_6
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ replica_cell_1rw
Xrbc_7
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ replica_cell_1rw
Xrbc_8
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ replica_cell_1rw
Xrbc_9
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ replica_cell_1rw
Xrbc_10
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ replica_cell_1rw
Xrbc_11
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ replica_cell_1rw
Xrbc_12
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ replica_cell_1rw
Xrbc_13
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ replica_cell_1rw
Xrbc_14
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ replica_cell_1rw
Xrbc_15
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ replica_cell_1rw
Xrbc_16
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ replica_cell_1rw
Xrbc_17
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ replica_cell_1rw
Xrbc_18
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ replica_cell_1rw
Xrbc_19
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ replica_cell_1rw
Xrbc_20
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ replica_cell_1rw
Xrbc_21
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ replica_cell_1rw
Xrbc_22
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ replica_cell_1rw
Xrbc_23
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ replica_cell_1rw
Xrbc_24
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ replica_cell_1rw
Xrbc_25
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ replica_cell_1rw
Xrbc_26
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ replica_cell_1rw
Xrbc_27
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ replica_cell_1rw
Xrbc_28
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ replica_cell_1rw
Xrbc_29
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ replica_cell_1rw
Xrbc_30
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ replica_cell_1rw
Xrbc_31
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ replica_cell_1rw
Xrbc_32
+ bl_0_0 br_0_0 wl_0_32 vdd gnd
+ replica_cell_1rw
.ENDS scn4m_subm_256x8_replica_column

*********************** "cell_1rw" ******************************
.SUBCKT cell_1rw bl br wl vdd gnd
* SPICE3 file created from cell_1rw.ext - technology: scmos

* Inverter 1
M1000 Q Q_bar vdd vdd p w=0.6u l=0.8u
M1002 Q Q_bar gnd gnd n w=1.6u l=0.4u

* Inverter 2
M1001 vdd Q Q_bar vdd p w=0.6u l=0.8u
M1003 gnd Q Q_bar gnd n w=1.6u l=0.4u

* Access transistors
M1004 Q wl bl gnd n w=0.8u l=0.4u
M1005 Q_bar wl br gnd n w=0.8u l=0.4u

.ENDS

.SUBCKT scn4m_subm_256x8_bitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* POWER : vdd 
* GROUND: gnd 
* rows: 32 cols: 64
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c0
+ bl_0_0 br_0_0 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c0
+ bl_0_0 br_0_0 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c0
+ bl_0_0 br_0_0 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c0
+ bl_0_0 br_0_0 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c0
+ bl_0_0 br_0_0 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c0
+ bl_0_0 br_0_0 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c0
+ bl_0_0 br_0_0 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c0
+ bl_0_0 br_0_0 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c0
+ bl_0_0 br_0_0 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c0
+ bl_0_0 br_0_0 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c0
+ bl_0_0 br_0_0 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c0
+ bl_0_0 br_0_0 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c0
+ bl_0_0 br_0_0 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c0
+ bl_0_0 br_0_0 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c0
+ bl_0_0 br_0_0 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c0
+ bl_0_0 br_0_0 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c0
+ bl_0_0 br_0_0 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c0
+ bl_0_0 br_0_0 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c0
+ bl_0_0 br_0_0 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c0
+ bl_0_0 br_0_0 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c0
+ bl_0_0 br_0_0 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c0
+ bl_0_0 br_0_0 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c0
+ bl_0_0 br_0_0 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c0
+ bl_0_0 br_0_0 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c0
+ bl_0_0 br_0_0 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c0
+ bl_0_0 br_0_0 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c0
+ bl_0_0 br_0_0 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c0
+ bl_0_0 br_0_0 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c0
+ bl_0_0 br_0_0 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c0
+ bl_0_0 br_0_0 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c0
+ bl_0_0 br_0_0 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c1
*+ bl_0_1 br_0_1 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c1
*+ bl_0_1 br_0_1 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c1
*+ bl_0_1 br_0_1 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c1
*+ bl_0_1 br_0_1 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c1
*+ bl_0_1 br_0_1 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c1
*+ bl_0_1 br_0_1 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c1
*+ bl_0_1 br_0_1 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c1
*+ bl_0_1 br_0_1 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c1
*+ bl_0_1 br_0_1 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c1
*+ bl_0_1 br_0_1 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c1
*+ bl_0_1 br_0_1 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c1
*+ bl_0_1 br_0_1 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c1
*+ bl_0_1 br_0_1 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c1
*+ bl_0_1 br_0_1 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c1
*+ bl_0_1 br_0_1 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c1
*+ bl_0_1 br_0_1 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c1
*+ bl_0_1 br_0_1 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c1
*+ bl_0_1 br_0_1 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c1
*+ bl_0_1 br_0_1 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c1
*+ bl_0_1 br_0_1 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c1
*+ bl_0_1 br_0_1 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c1
*+ bl_0_1 br_0_1 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c1
*+ bl_0_1 br_0_1 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c1
*+ bl_0_1 br_0_1 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c1
*+ bl_0_1 br_0_1 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c1
*+ bl_0_1 br_0_1 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c1
*+ bl_0_1 br_0_1 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c1
*+ bl_0_1 br_0_1 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c1
*+ bl_0_1 br_0_1 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c1
*+ bl_0_1 br_0_1 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c1
+ bl_0_1 br_0_1 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c2
*+ bl_0_2 br_0_2 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c2
*+ bl_0_2 br_0_2 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c2
*+ bl_0_2 br_0_2 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c2
*+ bl_0_2 br_0_2 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c2
*+ bl_0_2 br_0_2 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c2
*+ bl_0_2 br_0_2 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c2
*+ bl_0_2 br_0_2 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c2
*+ bl_0_2 br_0_2 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c2
*+ bl_0_2 br_0_2 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c2
*+ bl_0_2 br_0_2 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c2
*+ bl_0_2 br_0_2 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c2
*+ bl_0_2 br_0_2 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c2
*+ bl_0_2 br_0_2 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c2
*+ bl_0_2 br_0_2 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c2
*+ bl_0_2 br_0_2 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c2
*+ bl_0_2 br_0_2 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c2
*+ bl_0_2 br_0_2 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c2
*+ bl_0_2 br_0_2 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c2
*+ bl_0_2 br_0_2 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c2
*+ bl_0_2 br_0_2 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c2
*+ bl_0_2 br_0_2 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c2
*+ bl_0_2 br_0_2 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c2
*+ bl_0_2 br_0_2 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c2
*+ bl_0_2 br_0_2 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c2
*+ bl_0_2 br_0_2 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c2
*+ bl_0_2 br_0_2 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c2
*+ bl_0_2 br_0_2 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c2
*+ bl_0_2 br_0_2 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c2
*+ bl_0_2 br_0_2 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c2
*+ bl_0_2 br_0_2 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c2
+ bl_0_2 br_0_2 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c3
*+ bl_0_3 br_0_3 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c3
*+ bl_0_3 br_0_3 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c3
*+ bl_0_3 br_0_3 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c3
*+ bl_0_3 br_0_3 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c3
*+ bl_0_3 br_0_3 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c3
*+ bl_0_3 br_0_3 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c3
*+ bl_0_3 br_0_3 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c3
*+ bl_0_3 br_0_3 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c3
*+ bl_0_3 br_0_3 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c3
*+ bl_0_3 br_0_3 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c3
*+ bl_0_3 br_0_3 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c3
*+ bl_0_3 br_0_3 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c3
*+ bl_0_3 br_0_3 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c3
*+ bl_0_3 br_0_3 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c3
*+ bl_0_3 br_0_3 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c3
*+ bl_0_3 br_0_3 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c3
*+ bl_0_3 br_0_3 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c3
*+ bl_0_3 br_0_3 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c3
*+ bl_0_3 br_0_3 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c3
*+ bl_0_3 br_0_3 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c3
*+ bl_0_3 br_0_3 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c3
*+ bl_0_3 br_0_3 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c3
*+ bl_0_3 br_0_3 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c3
*+ bl_0_3 br_0_3 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c3
*+ bl_0_3 br_0_3 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c3
*+ bl_0_3 br_0_3 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c3
*+ bl_0_3 br_0_3 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c3
*+ bl_0_3 br_0_3 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c3
*+ bl_0_3 br_0_3 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c3
*+ bl_0_3 br_0_3 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c3
+ bl_0_3 br_0_3 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c4
*+ bl_0_4 br_0_4 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c4
*+ bl_0_4 br_0_4 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c4
*+ bl_0_4 br_0_4 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c4
*+ bl_0_4 br_0_4 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c4
*+ bl_0_4 br_0_4 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c4
*+ bl_0_4 br_0_4 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c4
*+ bl_0_4 br_0_4 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c4
*+ bl_0_4 br_0_4 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c4
*+ bl_0_4 br_0_4 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c4
*+ bl_0_4 br_0_4 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c4
*+ bl_0_4 br_0_4 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c4
*+ bl_0_4 br_0_4 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c4
*+ bl_0_4 br_0_4 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c4
*+ bl_0_4 br_0_4 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c4
*+ bl_0_4 br_0_4 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c4
*+ bl_0_4 br_0_4 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c4
*+ bl_0_4 br_0_4 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c4
*+ bl_0_4 br_0_4 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c4
*+ bl_0_4 br_0_4 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c4
*+ bl_0_4 br_0_4 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c4
*+ bl_0_4 br_0_4 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c4
*+ bl_0_4 br_0_4 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c4
*+ bl_0_4 br_0_4 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c4
*+ bl_0_4 br_0_4 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c4
*+ bl_0_4 br_0_4 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c4
*+ bl_0_4 br_0_4 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c4
*+ bl_0_4 br_0_4 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c4
*+ bl_0_4 br_0_4 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c4
*+ bl_0_4 br_0_4 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c4
*+ bl_0_4 br_0_4 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c4
+ bl_0_4 br_0_4 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c5
*+ bl_0_5 br_0_5 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c5
*+ bl_0_5 br_0_5 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c5
*+ bl_0_5 br_0_5 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c5
*+ bl_0_5 br_0_5 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c5
*+ bl_0_5 br_0_5 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c5
*+ bl_0_5 br_0_5 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c5
*+ bl_0_5 br_0_5 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c5
*+ bl_0_5 br_0_5 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c5
*+ bl_0_5 br_0_5 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c5
*+ bl_0_5 br_0_5 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c5
*+ bl_0_5 br_0_5 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c5
*+ bl_0_5 br_0_5 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c5
*+ bl_0_5 br_0_5 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c5
*+ bl_0_5 br_0_5 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c5
*+ bl_0_5 br_0_5 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c5
*+ bl_0_5 br_0_5 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c5
*+ bl_0_5 br_0_5 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c5
*+ bl_0_5 br_0_5 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c5
*+ bl_0_5 br_0_5 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c5
*+ bl_0_5 br_0_5 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c5
*+ bl_0_5 br_0_5 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c5
*+ bl_0_5 br_0_5 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c5
*+ bl_0_5 br_0_5 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c5
*+ bl_0_5 br_0_5 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c5
*+ bl_0_5 br_0_5 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c5
*+ bl_0_5 br_0_5 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c5
*+ bl_0_5 br_0_5 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c5
*+ bl_0_5 br_0_5 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c5
*+ bl_0_5 br_0_5 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c5
*+ bl_0_5 br_0_5 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c5
+ bl_0_5 br_0_5 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c6
*+ bl_0_6 br_0_6 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c6
*+ bl_0_6 br_0_6 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c6
*+ bl_0_6 br_0_6 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c6
*+ bl_0_6 br_0_6 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c6
*+ bl_0_6 br_0_6 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c6
*+ bl_0_6 br_0_6 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c6
*+ bl_0_6 br_0_6 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c6
*+ bl_0_6 br_0_6 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c6
*+ bl_0_6 br_0_6 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c6
*+ bl_0_6 br_0_6 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c6
*+ bl_0_6 br_0_6 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c6
*+ bl_0_6 br_0_6 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c6
*+ bl_0_6 br_0_6 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c6
*+ bl_0_6 br_0_6 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c6
*+ bl_0_6 br_0_6 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c6
*+ bl_0_6 br_0_6 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c6
*+ bl_0_6 br_0_6 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c6
*+ bl_0_6 br_0_6 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c6
*+ bl_0_6 br_0_6 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c6
*+ bl_0_6 br_0_6 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c6
*+ bl_0_6 br_0_6 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c6
*+ bl_0_6 br_0_6 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c6
*+ bl_0_6 br_0_6 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c6
*+ bl_0_6 br_0_6 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c6
*+ bl_0_6 br_0_6 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c6
*+ bl_0_6 br_0_6 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c6
*+ bl_0_6 br_0_6 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c6
*+ bl_0_6 br_0_6 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c6
*+ bl_0_6 br_0_6 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c6
*+ bl_0_6 br_0_6 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c6
+ bl_0_6 br_0_6 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c7
*+ bl_0_7 br_0_7 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c7
*+ bl_0_7 br_0_7 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c7
*+ bl_0_7 br_0_7 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c7
*+ bl_0_7 br_0_7 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c7
*+ bl_0_7 br_0_7 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c7
*+ bl_0_7 br_0_7 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c7
*+ bl_0_7 br_0_7 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c7
*+ bl_0_7 br_0_7 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c7
*+ bl_0_7 br_0_7 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c7
*+ bl_0_7 br_0_7 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c7
*+ bl_0_7 br_0_7 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c7
*+ bl_0_7 br_0_7 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c7
*+ bl_0_7 br_0_7 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c7
*+ bl_0_7 br_0_7 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c7
*+ bl_0_7 br_0_7 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c7
*+ bl_0_7 br_0_7 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c7
*+ bl_0_7 br_0_7 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c7
*+ bl_0_7 br_0_7 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c7
*+ bl_0_7 br_0_7 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c7
*+ bl_0_7 br_0_7 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c7
*+ bl_0_7 br_0_7 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c7
*+ bl_0_7 br_0_7 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c7
*+ bl_0_7 br_0_7 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c7
*+ bl_0_7 br_0_7 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c7
*+ bl_0_7 br_0_7 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c7
*+ bl_0_7 br_0_7 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c7
*+ bl_0_7 br_0_7 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c7
*+ bl_0_7 br_0_7 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c7
*+ bl_0_7 br_0_7 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c7
*+ bl_0_7 br_0_7 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c7
+ bl_0_7 br_0_7 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c8
*+ bl_0_8 br_0_8 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c8
*+ bl_0_8 br_0_8 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c8
*+ bl_0_8 br_0_8 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c8
*+ bl_0_8 br_0_8 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c8
*+ bl_0_8 br_0_8 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c8
*+ bl_0_8 br_0_8 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c8
*+ bl_0_8 br_0_8 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c8
*+ bl_0_8 br_0_8 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c8
*+ bl_0_8 br_0_8 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c8
*+ bl_0_8 br_0_8 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c8
*+ bl_0_8 br_0_8 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c8
*+ bl_0_8 br_0_8 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c8
*+ bl_0_8 br_0_8 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c8
*+ bl_0_8 br_0_8 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c8
*+ bl_0_8 br_0_8 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c8
*+ bl_0_8 br_0_8 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c8
*+ bl_0_8 br_0_8 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c8
*+ bl_0_8 br_0_8 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c8
*+ bl_0_8 br_0_8 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c8
*+ bl_0_8 br_0_8 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c8
*+ bl_0_8 br_0_8 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c8
*+ bl_0_8 br_0_8 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c8
*+ bl_0_8 br_0_8 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c8
*+ bl_0_8 br_0_8 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c8
*+ bl_0_8 br_0_8 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c8
*+ bl_0_8 br_0_8 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c8
*+ bl_0_8 br_0_8 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c8
*+ bl_0_8 br_0_8 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c8
*+ bl_0_8 br_0_8 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c8
*+ bl_0_8 br_0_8 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c8
+ bl_0_8 br_0_8 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c9
*+ bl_0_9 br_0_9 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c9
*+ bl_0_9 br_0_9 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c9
*+ bl_0_9 br_0_9 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c9
*+ bl_0_9 br_0_9 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c9
*+ bl_0_9 br_0_9 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c9
*+ bl_0_9 br_0_9 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c9
*+ bl_0_9 br_0_9 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c9
*+ bl_0_9 br_0_9 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c9
*+ bl_0_9 br_0_9 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c9
*+ bl_0_9 br_0_9 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c9
*+ bl_0_9 br_0_9 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c9
*+ bl_0_9 br_0_9 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c9
*+ bl_0_9 br_0_9 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c9
*+ bl_0_9 br_0_9 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c9
*+ bl_0_9 br_0_9 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c9
*+ bl_0_9 br_0_9 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c9
*+ bl_0_9 br_0_9 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c9
*+ bl_0_9 br_0_9 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c9
*+ bl_0_9 br_0_9 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c9
*+ bl_0_9 br_0_9 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c9
*+ bl_0_9 br_0_9 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c9
*+ bl_0_9 br_0_9 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c9
*+ bl_0_9 br_0_9 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c9
*+ bl_0_9 br_0_9 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c9
*+ bl_0_9 br_0_9 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c9
*+ bl_0_9 br_0_9 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c9
*+ bl_0_9 br_0_9 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c9
*+ bl_0_9 br_0_9 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c9
*+ bl_0_9 br_0_9 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c9
*+ bl_0_9 br_0_9 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c9
+ bl_0_9 br_0_9 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c10
*+ bl_0_10 br_0_10 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c10
*+ bl_0_10 br_0_10 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c10
*+ bl_0_10 br_0_10 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c10
*+ bl_0_10 br_0_10 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c10
*+ bl_0_10 br_0_10 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c10
*+ bl_0_10 br_0_10 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c10
*+ bl_0_10 br_0_10 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c10
*+ bl_0_10 br_0_10 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c10
*+ bl_0_10 br_0_10 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c10
*+ bl_0_10 br_0_10 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c10
*+ bl_0_10 br_0_10 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c10
*+ bl_0_10 br_0_10 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c10
*+ bl_0_10 br_0_10 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c10
*+ bl_0_10 br_0_10 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c10
*+ bl_0_10 br_0_10 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c10
*+ bl_0_10 br_0_10 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c10
*+ bl_0_10 br_0_10 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c10
*+ bl_0_10 br_0_10 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c10
*+ bl_0_10 br_0_10 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c10
*+ bl_0_10 br_0_10 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c10
*+ bl_0_10 br_0_10 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c10
*+ bl_0_10 br_0_10 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c10
*+ bl_0_10 br_0_10 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c10
*+ bl_0_10 br_0_10 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c10
*+ bl_0_10 br_0_10 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c10
*+ bl_0_10 br_0_10 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c10
*+ bl_0_10 br_0_10 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c10
*+ bl_0_10 br_0_10 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c10
*+ bl_0_10 br_0_10 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c10
*+ bl_0_10 br_0_10 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c10
+ bl_0_10 br_0_10 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c11
*+ bl_0_11 br_0_11 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c11
*+ bl_0_11 br_0_11 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c11
*+ bl_0_11 br_0_11 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c11
*+ bl_0_11 br_0_11 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c11
*+ bl_0_11 br_0_11 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c11
*+ bl_0_11 br_0_11 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c11
*+ bl_0_11 br_0_11 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c11
*+ bl_0_11 br_0_11 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c11
*+ bl_0_11 br_0_11 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c11
*+ bl_0_11 br_0_11 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c11
*+ bl_0_11 br_0_11 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c11
*+ bl_0_11 br_0_11 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c11
*+ bl_0_11 br_0_11 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c11
*+ bl_0_11 br_0_11 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c11
*+ bl_0_11 br_0_11 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c11
*+ bl_0_11 br_0_11 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c11
*+ bl_0_11 br_0_11 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c11
*+ bl_0_11 br_0_11 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c11
*+ bl_0_11 br_0_11 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c11
*+ bl_0_11 br_0_11 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c11
*+ bl_0_11 br_0_11 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c11
*+ bl_0_11 br_0_11 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c11
*+ bl_0_11 br_0_11 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c11
*+ bl_0_11 br_0_11 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c11
*+ bl_0_11 br_0_11 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c11
*+ bl_0_11 br_0_11 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c11
*+ bl_0_11 br_0_11 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c11
*+ bl_0_11 br_0_11 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c11
*+ bl_0_11 br_0_11 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c11
*+ bl_0_11 br_0_11 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c11
+ bl_0_11 br_0_11 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c12
*+ bl_0_12 br_0_12 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c12
*+ bl_0_12 br_0_12 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c12
*+ bl_0_12 br_0_12 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c12
*+ bl_0_12 br_0_12 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c12
*+ bl_0_12 br_0_12 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c12
*+ bl_0_12 br_0_12 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c12
*+ bl_0_12 br_0_12 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c12
*+ bl_0_12 br_0_12 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c12
*+ bl_0_12 br_0_12 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c12
*+ bl_0_12 br_0_12 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c12
*+ bl_0_12 br_0_12 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c12
*+ bl_0_12 br_0_12 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c12
*+ bl_0_12 br_0_12 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c12
*+ bl_0_12 br_0_12 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c12
*+ bl_0_12 br_0_12 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c12
*+ bl_0_12 br_0_12 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c12
*+ bl_0_12 br_0_12 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c12
*+ bl_0_12 br_0_12 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c12
*+ bl_0_12 br_0_12 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c12
*+ bl_0_12 br_0_12 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c12
*+ bl_0_12 br_0_12 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c12
*+ bl_0_12 br_0_12 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c12
*+ bl_0_12 br_0_12 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c12
*+ bl_0_12 br_0_12 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c12
*+ bl_0_12 br_0_12 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c12
*+ bl_0_12 br_0_12 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c12
*+ bl_0_12 br_0_12 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c12
*+ bl_0_12 br_0_12 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c12
*+ bl_0_12 br_0_12 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c12
*+ bl_0_12 br_0_12 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c12
+ bl_0_12 br_0_12 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c13
*+ bl_0_13 br_0_13 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c13
*+ bl_0_13 br_0_13 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c13
*+ bl_0_13 br_0_13 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c13
*+ bl_0_13 br_0_13 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c13
*+ bl_0_13 br_0_13 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c13
*+ bl_0_13 br_0_13 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c13
*+ bl_0_13 br_0_13 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c13
*+ bl_0_13 br_0_13 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c13
*+ bl_0_13 br_0_13 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c13
*+ bl_0_13 br_0_13 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c13
*+ bl_0_13 br_0_13 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c13
*+ bl_0_13 br_0_13 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c13
*+ bl_0_13 br_0_13 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c13
*+ bl_0_13 br_0_13 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c13
*+ bl_0_13 br_0_13 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c13
*+ bl_0_13 br_0_13 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c13
*+ bl_0_13 br_0_13 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c13
*+ bl_0_13 br_0_13 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c13
*+ bl_0_13 br_0_13 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c13
*+ bl_0_13 br_0_13 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c13
*+ bl_0_13 br_0_13 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c13
*+ bl_0_13 br_0_13 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c13
*+ bl_0_13 br_0_13 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c13
*+ bl_0_13 br_0_13 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c13
*+ bl_0_13 br_0_13 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c13
*+ bl_0_13 br_0_13 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c13
*+ bl_0_13 br_0_13 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c13
*+ bl_0_13 br_0_13 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c13
*+ bl_0_13 br_0_13 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c13
*+ bl_0_13 br_0_13 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c13
+ bl_0_13 br_0_13 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c14
*+ bl_0_14 br_0_14 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c14
*+ bl_0_14 br_0_14 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c14
*+ bl_0_14 br_0_14 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c14
*+ bl_0_14 br_0_14 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c14
*+ bl_0_14 br_0_14 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c14
*+ bl_0_14 br_0_14 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c14
*+ bl_0_14 br_0_14 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c14
*+ bl_0_14 br_0_14 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c14
*+ bl_0_14 br_0_14 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c14
*+ bl_0_14 br_0_14 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c14
*+ bl_0_14 br_0_14 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c14
*+ bl_0_14 br_0_14 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c14
*+ bl_0_14 br_0_14 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c14
*+ bl_0_14 br_0_14 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c14
*+ bl_0_14 br_0_14 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c14
*+ bl_0_14 br_0_14 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c14
*+ bl_0_14 br_0_14 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c14
*+ bl_0_14 br_0_14 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c14
*+ bl_0_14 br_0_14 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c14
*+ bl_0_14 br_0_14 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c14
*+ bl_0_14 br_0_14 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c14
*+ bl_0_14 br_0_14 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c14
*+ bl_0_14 br_0_14 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c14
*+ bl_0_14 br_0_14 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c14
*+ bl_0_14 br_0_14 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c14
*+ bl_0_14 br_0_14 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c14
*+ bl_0_14 br_0_14 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c14
*+ bl_0_14 br_0_14 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c14
*+ bl_0_14 br_0_14 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c14
*+ bl_0_14 br_0_14 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c14
+ bl_0_14 br_0_14 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c15
*+ bl_0_15 br_0_15 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c15
*+ bl_0_15 br_0_15 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c15
*+ bl_0_15 br_0_15 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c15
*+ bl_0_15 br_0_15 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c15
*+ bl_0_15 br_0_15 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c15
*+ bl_0_15 br_0_15 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c15
*+ bl_0_15 br_0_15 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c15
*+ bl_0_15 br_0_15 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c15
*+ bl_0_15 br_0_15 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c15
*+ bl_0_15 br_0_15 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c15
*+ bl_0_15 br_0_15 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c15
*+ bl_0_15 br_0_15 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c15
*+ bl_0_15 br_0_15 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c15
*+ bl_0_15 br_0_15 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c15
*+ bl_0_15 br_0_15 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c15
*+ bl_0_15 br_0_15 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c15
*+ bl_0_15 br_0_15 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c15
*+ bl_0_15 br_0_15 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c15
*+ bl_0_15 br_0_15 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c15
*+ bl_0_15 br_0_15 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c15
*+ bl_0_15 br_0_15 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c15
*+ bl_0_15 br_0_15 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c15
*+ bl_0_15 br_0_15 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c15
*+ bl_0_15 br_0_15 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c15
*+ bl_0_15 br_0_15 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c15
*+ bl_0_15 br_0_15 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c15
*+ bl_0_15 br_0_15 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c15
*+ bl_0_15 br_0_15 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c15
*+ bl_0_15 br_0_15 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c15
*+ bl_0_15 br_0_15 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c15
+ bl_0_15 br_0_15 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c16
*+ bl_0_16 br_0_16 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c16
*+ bl_0_16 br_0_16 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c16
*+ bl_0_16 br_0_16 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c16
*+ bl_0_16 br_0_16 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c16
*+ bl_0_16 br_0_16 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c16
*+ bl_0_16 br_0_16 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c16
*+ bl_0_16 br_0_16 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c16
*+ bl_0_16 br_0_16 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c16
*+ bl_0_16 br_0_16 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c16
*+ bl_0_16 br_0_16 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c16
*+ bl_0_16 br_0_16 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c16
*+ bl_0_16 br_0_16 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c16
*+ bl_0_16 br_0_16 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c16
*+ bl_0_16 br_0_16 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c16
*+ bl_0_16 br_0_16 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c16
*+ bl_0_16 br_0_16 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c16
*+ bl_0_16 br_0_16 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c16
*+ bl_0_16 br_0_16 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c16
*+ bl_0_16 br_0_16 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c16
*+ bl_0_16 br_0_16 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c16
*+ bl_0_16 br_0_16 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c16
*+ bl_0_16 br_0_16 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c16
*+ bl_0_16 br_0_16 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c16
*+ bl_0_16 br_0_16 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c16
*+ bl_0_16 br_0_16 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c16
*+ bl_0_16 br_0_16 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c16
*+ bl_0_16 br_0_16 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c16
*+ bl_0_16 br_0_16 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c16
*+ bl_0_16 br_0_16 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c16
*+ bl_0_16 br_0_16 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c16
+ bl_0_16 br_0_16 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c17
*+ bl_0_17 br_0_17 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c17
*+ bl_0_17 br_0_17 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c17
*+ bl_0_17 br_0_17 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c17
*+ bl_0_17 br_0_17 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c17
*+ bl_0_17 br_0_17 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c17
*+ bl_0_17 br_0_17 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c17
*+ bl_0_17 br_0_17 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c17
*+ bl_0_17 br_0_17 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c17
*+ bl_0_17 br_0_17 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c17
*+ bl_0_17 br_0_17 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c17
*+ bl_0_17 br_0_17 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c17
*+ bl_0_17 br_0_17 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c17
*+ bl_0_17 br_0_17 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c17
*+ bl_0_17 br_0_17 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c17
*+ bl_0_17 br_0_17 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c17
*+ bl_0_17 br_0_17 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c17
*+ bl_0_17 br_0_17 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c17
*+ bl_0_17 br_0_17 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c17
*+ bl_0_17 br_0_17 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c17
*+ bl_0_17 br_0_17 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c17
*+ bl_0_17 br_0_17 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c17
*+ bl_0_17 br_0_17 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c17
*+ bl_0_17 br_0_17 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c17
*+ bl_0_17 br_0_17 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c17
*+ bl_0_17 br_0_17 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c17
*+ bl_0_17 br_0_17 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c17
*+ bl_0_17 br_0_17 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c17
*+ bl_0_17 br_0_17 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c17
*+ bl_0_17 br_0_17 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c17
*+ bl_0_17 br_0_17 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c17
+ bl_0_17 br_0_17 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c18
*+ bl_0_18 br_0_18 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c18
*+ bl_0_18 br_0_18 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c18
*+ bl_0_18 br_0_18 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c18
*+ bl_0_18 br_0_18 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c18
*+ bl_0_18 br_0_18 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c18
*+ bl_0_18 br_0_18 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c18
*+ bl_0_18 br_0_18 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c18
*+ bl_0_18 br_0_18 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c18
*+ bl_0_18 br_0_18 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c18
*+ bl_0_18 br_0_18 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c18
*+ bl_0_18 br_0_18 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c18
*+ bl_0_18 br_0_18 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c18
*+ bl_0_18 br_0_18 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c18
*+ bl_0_18 br_0_18 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c18
*+ bl_0_18 br_0_18 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c18
*+ bl_0_18 br_0_18 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c18
*+ bl_0_18 br_0_18 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c18
*+ bl_0_18 br_0_18 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c18
*+ bl_0_18 br_0_18 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c18
*+ bl_0_18 br_0_18 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c18
*+ bl_0_18 br_0_18 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c18
*+ bl_0_18 br_0_18 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c18
*+ bl_0_18 br_0_18 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c18
*+ bl_0_18 br_0_18 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c18
*+ bl_0_18 br_0_18 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c18
*+ bl_0_18 br_0_18 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c18
*+ bl_0_18 br_0_18 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c18
*+ bl_0_18 br_0_18 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c18
*+ bl_0_18 br_0_18 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c18
*+ bl_0_18 br_0_18 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c18
+ bl_0_18 br_0_18 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c19
*+ bl_0_19 br_0_19 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c19
*+ bl_0_19 br_0_19 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c19
*+ bl_0_19 br_0_19 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c19
*+ bl_0_19 br_0_19 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c19
*+ bl_0_19 br_0_19 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c19
*+ bl_0_19 br_0_19 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c19
*+ bl_0_19 br_0_19 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c19
*+ bl_0_19 br_0_19 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c19
*+ bl_0_19 br_0_19 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c19
*+ bl_0_19 br_0_19 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c19
*+ bl_0_19 br_0_19 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c19
*+ bl_0_19 br_0_19 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c19
*+ bl_0_19 br_0_19 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c19
*+ bl_0_19 br_0_19 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c19
*+ bl_0_19 br_0_19 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c19
*+ bl_0_19 br_0_19 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c19
*+ bl_0_19 br_0_19 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c19
*+ bl_0_19 br_0_19 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c19
*+ bl_0_19 br_0_19 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c19
*+ bl_0_19 br_0_19 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c19
*+ bl_0_19 br_0_19 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c19
*+ bl_0_19 br_0_19 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c19
*+ bl_0_19 br_0_19 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c19
*+ bl_0_19 br_0_19 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c19
*+ bl_0_19 br_0_19 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c19
*+ bl_0_19 br_0_19 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c19
*+ bl_0_19 br_0_19 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c19
*+ bl_0_19 br_0_19 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c19
*+ bl_0_19 br_0_19 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c19
*+ bl_0_19 br_0_19 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c19
+ bl_0_19 br_0_19 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c20
*+ bl_0_20 br_0_20 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c20
*+ bl_0_20 br_0_20 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c20
*+ bl_0_20 br_0_20 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c20
*+ bl_0_20 br_0_20 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c20
*+ bl_0_20 br_0_20 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c20
*+ bl_0_20 br_0_20 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c20
*+ bl_0_20 br_0_20 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c20
*+ bl_0_20 br_0_20 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c20
*+ bl_0_20 br_0_20 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c20
*+ bl_0_20 br_0_20 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c20
*+ bl_0_20 br_0_20 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c20
*+ bl_0_20 br_0_20 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c20
*+ bl_0_20 br_0_20 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c20
*+ bl_0_20 br_0_20 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c20
*+ bl_0_20 br_0_20 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c20
*+ bl_0_20 br_0_20 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c20
*+ bl_0_20 br_0_20 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c20
*+ bl_0_20 br_0_20 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c20
*+ bl_0_20 br_0_20 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c20
*+ bl_0_20 br_0_20 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c20
*+ bl_0_20 br_0_20 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c20
*+ bl_0_20 br_0_20 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c20
*+ bl_0_20 br_0_20 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c20
*+ bl_0_20 br_0_20 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c20
*+ bl_0_20 br_0_20 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c20
*+ bl_0_20 br_0_20 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c20
*+ bl_0_20 br_0_20 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c20
*+ bl_0_20 br_0_20 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c20
*+ bl_0_20 br_0_20 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c20
*+ bl_0_20 br_0_20 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c20
+ bl_0_20 br_0_20 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c21
*+ bl_0_21 br_0_21 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c21
*+ bl_0_21 br_0_21 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c21
*+ bl_0_21 br_0_21 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c21
*+ bl_0_21 br_0_21 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c21
*+ bl_0_21 br_0_21 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c21
*+ bl_0_21 br_0_21 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c21
*+ bl_0_21 br_0_21 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c21
*+ bl_0_21 br_0_21 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c21
*+ bl_0_21 br_0_21 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c21
*+ bl_0_21 br_0_21 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c21
*+ bl_0_21 br_0_21 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c21
*+ bl_0_21 br_0_21 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c21
*+ bl_0_21 br_0_21 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c21
*+ bl_0_21 br_0_21 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c21
*+ bl_0_21 br_0_21 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c21
*+ bl_0_21 br_0_21 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c21
*+ bl_0_21 br_0_21 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c21
*+ bl_0_21 br_0_21 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c21
*+ bl_0_21 br_0_21 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c21
*+ bl_0_21 br_0_21 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c21
*+ bl_0_21 br_0_21 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c21
*+ bl_0_21 br_0_21 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c21
*+ bl_0_21 br_0_21 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c21
*+ bl_0_21 br_0_21 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c21
*+ bl_0_21 br_0_21 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c21
*+ bl_0_21 br_0_21 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c21
*+ bl_0_21 br_0_21 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c21
*+ bl_0_21 br_0_21 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c21
*+ bl_0_21 br_0_21 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c21
*+ bl_0_21 br_0_21 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c21
+ bl_0_21 br_0_21 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c22
*+ bl_0_22 br_0_22 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c22
*+ bl_0_22 br_0_22 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c22
*+ bl_0_22 br_0_22 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c22
*+ bl_0_22 br_0_22 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c22
*+ bl_0_22 br_0_22 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c22
*+ bl_0_22 br_0_22 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c22
*+ bl_0_22 br_0_22 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c22
*+ bl_0_22 br_0_22 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c22
*+ bl_0_22 br_0_22 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c22
*+ bl_0_22 br_0_22 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c22
*+ bl_0_22 br_0_22 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c22
*+ bl_0_22 br_0_22 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c22
*+ bl_0_22 br_0_22 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c22
*+ bl_0_22 br_0_22 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c22
*+ bl_0_22 br_0_22 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c22
*+ bl_0_22 br_0_22 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c22
*+ bl_0_22 br_0_22 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c22
*+ bl_0_22 br_0_22 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c22
*+ bl_0_22 br_0_22 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c22
*+ bl_0_22 br_0_22 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c22
*+ bl_0_22 br_0_22 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c22
*+ bl_0_22 br_0_22 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c22
*+ bl_0_22 br_0_22 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c22
*+ bl_0_22 br_0_22 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c22
*+ bl_0_22 br_0_22 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c22
*+ bl_0_22 br_0_22 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c22
*+ bl_0_22 br_0_22 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c22
*+ bl_0_22 br_0_22 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c22
*+ bl_0_22 br_0_22 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c22
*+ bl_0_22 br_0_22 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c22
+ bl_0_22 br_0_22 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c23
*+ bl_0_23 br_0_23 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c23
*+ bl_0_23 br_0_23 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c23
*+ bl_0_23 br_0_23 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c23
*+ bl_0_23 br_0_23 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c23
*+ bl_0_23 br_0_23 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c23
*+ bl_0_23 br_0_23 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c23
*+ bl_0_23 br_0_23 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c23
*+ bl_0_23 br_0_23 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c23
*+ bl_0_23 br_0_23 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c23
*+ bl_0_23 br_0_23 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c23
*+ bl_0_23 br_0_23 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c23
*+ bl_0_23 br_0_23 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c23
*+ bl_0_23 br_0_23 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c23
*+ bl_0_23 br_0_23 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c23
*+ bl_0_23 br_0_23 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c23
*+ bl_0_23 br_0_23 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c23
*+ bl_0_23 br_0_23 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c23
*+ bl_0_23 br_0_23 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c23
*+ bl_0_23 br_0_23 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c23
*+ bl_0_23 br_0_23 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c23
*+ bl_0_23 br_0_23 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c23
*+ bl_0_23 br_0_23 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c23
*+ bl_0_23 br_0_23 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c23
*+ bl_0_23 br_0_23 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c23
*+ bl_0_23 br_0_23 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c23
*+ bl_0_23 br_0_23 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c23
*+ bl_0_23 br_0_23 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c23
*+ bl_0_23 br_0_23 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c23
*+ bl_0_23 br_0_23 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c23
*+ bl_0_23 br_0_23 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c23
+ bl_0_23 br_0_23 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c24
*+ bl_0_24 br_0_24 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c24
*+ bl_0_24 br_0_24 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c24
*+ bl_0_24 br_0_24 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c24
*+ bl_0_24 br_0_24 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c24
*+ bl_0_24 br_0_24 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c24
*+ bl_0_24 br_0_24 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c24
*+ bl_0_24 br_0_24 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c24
*+ bl_0_24 br_0_24 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c24
*+ bl_0_24 br_0_24 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c24
*+ bl_0_24 br_0_24 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c24
*+ bl_0_24 br_0_24 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c24
*+ bl_0_24 br_0_24 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c24
*+ bl_0_24 br_0_24 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c24
*+ bl_0_24 br_0_24 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c24
*+ bl_0_24 br_0_24 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c24
*+ bl_0_24 br_0_24 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c24
*+ bl_0_24 br_0_24 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c24
*+ bl_0_24 br_0_24 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c24
*+ bl_0_24 br_0_24 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c24
*+ bl_0_24 br_0_24 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c24
*+ bl_0_24 br_0_24 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c24
*+ bl_0_24 br_0_24 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c24
*+ bl_0_24 br_0_24 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c24
*+ bl_0_24 br_0_24 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c24
*+ bl_0_24 br_0_24 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c24
*+ bl_0_24 br_0_24 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c24
*+ bl_0_24 br_0_24 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c24
*+ bl_0_24 br_0_24 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c24
*+ bl_0_24 br_0_24 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c24
*+ bl_0_24 br_0_24 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c24
+ bl_0_24 br_0_24 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c25
*+ bl_0_25 br_0_25 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c25
*+ bl_0_25 br_0_25 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c25
*+ bl_0_25 br_0_25 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c25
*+ bl_0_25 br_0_25 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c25
*+ bl_0_25 br_0_25 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c25
*+ bl_0_25 br_0_25 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c25
*+ bl_0_25 br_0_25 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c25
*+ bl_0_25 br_0_25 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c25
*+ bl_0_25 br_0_25 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c25
*+ bl_0_25 br_0_25 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c25
*+ bl_0_25 br_0_25 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c25
*+ bl_0_25 br_0_25 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c25
*+ bl_0_25 br_0_25 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c25
*+ bl_0_25 br_0_25 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c25
*+ bl_0_25 br_0_25 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c25
*+ bl_0_25 br_0_25 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c25
*+ bl_0_25 br_0_25 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c25
*+ bl_0_25 br_0_25 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c25
*+ bl_0_25 br_0_25 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c25
*+ bl_0_25 br_0_25 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c25
*+ bl_0_25 br_0_25 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c25
*+ bl_0_25 br_0_25 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c25
*+ bl_0_25 br_0_25 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c25
*+ bl_0_25 br_0_25 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c25
*+ bl_0_25 br_0_25 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c25
*+ bl_0_25 br_0_25 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c25
*+ bl_0_25 br_0_25 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c25
*+ bl_0_25 br_0_25 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c25
*+ bl_0_25 br_0_25 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c25
*+ bl_0_25 br_0_25 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c25
+ bl_0_25 br_0_25 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c26
*+ bl_0_26 br_0_26 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c26
*+ bl_0_26 br_0_26 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c26
*+ bl_0_26 br_0_26 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c26
*+ bl_0_26 br_0_26 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c26
*+ bl_0_26 br_0_26 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c26
*+ bl_0_26 br_0_26 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c26
*+ bl_0_26 br_0_26 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c26
*+ bl_0_26 br_0_26 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c26
*+ bl_0_26 br_0_26 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c26
*+ bl_0_26 br_0_26 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c26
*+ bl_0_26 br_0_26 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c26
*+ bl_0_26 br_0_26 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c26
*+ bl_0_26 br_0_26 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c26
*+ bl_0_26 br_0_26 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c26
*+ bl_0_26 br_0_26 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c26
*+ bl_0_26 br_0_26 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c26
*+ bl_0_26 br_0_26 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c26
*+ bl_0_26 br_0_26 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c26
*+ bl_0_26 br_0_26 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c26
*+ bl_0_26 br_0_26 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c26
*+ bl_0_26 br_0_26 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c26
*+ bl_0_26 br_0_26 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c26
*+ bl_0_26 br_0_26 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c26
*+ bl_0_26 br_0_26 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c26
*+ bl_0_26 br_0_26 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c26
*+ bl_0_26 br_0_26 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c26
*+ bl_0_26 br_0_26 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c26
*+ bl_0_26 br_0_26 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c26
*+ bl_0_26 br_0_26 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c26
*+ bl_0_26 br_0_26 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c26
+ bl_0_26 br_0_26 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c27
*+ bl_0_27 br_0_27 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c27
*+ bl_0_27 br_0_27 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c27
*+ bl_0_27 br_0_27 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c27
*+ bl_0_27 br_0_27 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c27
*+ bl_0_27 br_0_27 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c27
*+ bl_0_27 br_0_27 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c27
*+ bl_0_27 br_0_27 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c27
*+ bl_0_27 br_0_27 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c27
*+ bl_0_27 br_0_27 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c27
*+ bl_0_27 br_0_27 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c27
*+ bl_0_27 br_0_27 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c27
*+ bl_0_27 br_0_27 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c27
*+ bl_0_27 br_0_27 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c27
*+ bl_0_27 br_0_27 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c27
*+ bl_0_27 br_0_27 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c27
*+ bl_0_27 br_0_27 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c27
*+ bl_0_27 br_0_27 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c27
*+ bl_0_27 br_0_27 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c27
*+ bl_0_27 br_0_27 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c27
*+ bl_0_27 br_0_27 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c27
*+ bl_0_27 br_0_27 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c27
*+ bl_0_27 br_0_27 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c27
*+ bl_0_27 br_0_27 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c27
*+ bl_0_27 br_0_27 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c27
*+ bl_0_27 br_0_27 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c27
*+ bl_0_27 br_0_27 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c27
*+ bl_0_27 br_0_27 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c27
*+ bl_0_27 br_0_27 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c27
*+ bl_0_27 br_0_27 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c27
*+ bl_0_27 br_0_27 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c27
+ bl_0_27 br_0_27 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c28
*+ bl_0_28 br_0_28 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c28
*+ bl_0_28 br_0_28 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c28
*+ bl_0_28 br_0_28 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c28
*+ bl_0_28 br_0_28 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c28
*+ bl_0_28 br_0_28 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c28
*+ bl_0_28 br_0_28 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c28
*+ bl_0_28 br_0_28 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c28
*+ bl_0_28 br_0_28 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c28
*+ bl_0_28 br_0_28 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c28
*+ bl_0_28 br_0_28 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c28
*+ bl_0_28 br_0_28 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c28
*+ bl_0_28 br_0_28 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c28
*+ bl_0_28 br_0_28 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c28
*+ bl_0_28 br_0_28 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c28
*+ bl_0_28 br_0_28 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c28
*+ bl_0_28 br_0_28 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c28
*+ bl_0_28 br_0_28 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c28
*+ bl_0_28 br_0_28 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c28
*+ bl_0_28 br_0_28 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c28
*+ bl_0_28 br_0_28 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c28
*+ bl_0_28 br_0_28 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c28
*+ bl_0_28 br_0_28 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c28
*+ bl_0_28 br_0_28 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c28
*+ bl_0_28 br_0_28 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c28
*+ bl_0_28 br_0_28 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c28
*+ bl_0_28 br_0_28 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c28
*+ bl_0_28 br_0_28 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c28
*+ bl_0_28 br_0_28 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c28
*+ bl_0_28 br_0_28 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c28
*+ bl_0_28 br_0_28 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c28
+ bl_0_28 br_0_28 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c29
*+ bl_0_29 br_0_29 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c29
*+ bl_0_29 br_0_29 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c29
*+ bl_0_29 br_0_29 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c29
*+ bl_0_29 br_0_29 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c29
*+ bl_0_29 br_0_29 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c29
*+ bl_0_29 br_0_29 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c29
*+ bl_0_29 br_0_29 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c29
*+ bl_0_29 br_0_29 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c29
*+ bl_0_29 br_0_29 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c29
*+ bl_0_29 br_0_29 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c29
*+ bl_0_29 br_0_29 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c29
*+ bl_0_29 br_0_29 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c29
*+ bl_0_29 br_0_29 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c29
*+ bl_0_29 br_0_29 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c29
*+ bl_0_29 br_0_29 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c29
*+ bl_0_29 br_0_29 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c29
*+ bl_0_29 br_0_29 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c29
*+ bl_0_29 br_0_29 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c29
*+ bl_0_29 br_0_29 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c29
*+ bl_0_29 br_0_29 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c29
*+ bl_0_29 br_0_29 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c29
*+ bl_0_29 br_0_29 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c29
*+ bl_0_29 br_0_29 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c29
*+ bl_0_29 br_0_29 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c29
*+ bl_0_29 br_0_29 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c29
*+ bl_0_29 br_0_29 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c29
*+ bl_0_29 br_0_29 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c29
*+ bl_0_29 br_0_29 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c29
*+ bl_0_29 br_0_29 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c29
*+ bl_0_29 br_0_29 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c29
+ bl_0_29 br_0_29 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c30
*+ bl_0_30 br_0_30 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c30
*+ bl_0_30 br_0_30 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c30
*+ bl_0_30 br_0_30 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c30
*+ bl_0_30 br_0_30 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c30
*+ bl_0_30 br_0_30 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c30
*+ bl_0_30 br_0_30 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c30
*+ bl_0_30 br_0_30 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c30
*+ bl_0_30 br_0_30 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c30
*+ bl_0_30 br_0_30 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c30
*+ bl_0_30 br_0_30 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c30
*+ bl_0_30 br_0_30 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c30
*+ bl_0_30 br_0_30 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c30
*+ bl_0_30 br_0_30 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c30
*+ bl_0_30 br_0_30 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c30
*+ bl_0_30 br_0_30 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c30
*+ bl_0_30 br_0_30 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c30
*+ bl_0_30 br_0_30 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c30
*+ bl_0_30 br_0_30 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c30
*+ bl_0_30 br_0_30 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c30
*+ bl_0_30 br_0_30 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c30
*+ bl_0_30 br_0_30 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c30
*+ bl_0_30 br_0_30 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c30
*+ bl_0_30 br_0_30 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c30
*+ bl_0_30 br_0_30 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c30
*+ bl_0_30 br_0_30 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c30
*+ bl_0_30 br_0_30 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c30
*+ bl_0_30 br_0_30 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c30
*+ bl_0_30 br_0_30 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c30
*+ bl_0_30 br_0_30 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c30
*+ bl_0_30 br_0_30 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c30
+ bl_0_30 br_0_30 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c31
*+ bl_0_31 br_0_31 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c31
*+ bl_0_31 br_0_31 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c31
*+ bl_0_31 br_0_31 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c31
*+ bl_0_31 br_0_31 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c31
*+ bl_0_31 br_0_31 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c31
*+ bl_0_31 br_0_31 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c31
*+ bl_0_31 br_0_31 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c31
*+ bl_0_31 br_0_31 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c31
*+ bl_0_31 br_0_31 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c31
*+ bl_0_31 br_0_31 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c31
*+ bl_0_31 br_0_31 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c31
*+ bl_0_31 br_0_31 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c31
*+ bl_0_31 br_0_31 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c31
*+ bl_0_31 br_0_31 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c31
*+ bl_0_31 br_0_31 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c31
*+ bl_0_31 br_0_31 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c31
*+ bl_0_31 br_0_31 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c31
*+ bl_0_31 br_0_31 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c31
*+ bl_0_31 br_0_31 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c31
*+ bl_0_31 br_0_31 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c31
*+ bl_0_31 br_0_31 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c31
*+ bl_0_31 br_0_31 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c31
*+ bl_0_31 br_0_31 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c31
*+ bl_0_31 br_0_31 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c31
*+ bl_0_31 br_0_31 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c31
*+ bl_0_31 br_0_31 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c31
*+ bl_0_31 br_0_31 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c31
*+ bl_0_31 br_0_31 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c31
*+ bl_0_31 br_0_31 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c31
*+ bl_0_31 br_0_31 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c31
+ bl_0_31 br_0_31 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c32
*+ bl_0_32 br_0_32 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c32
*+ bl_0_32 br_0_32 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c32
*+ bl_0_32 br_0_32 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c32
*+ bl_0_32 br_0_32 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c32
*+ bl_0_32 br_0_32 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c32
*+ bl_0_32 br_0_32 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c32
*+ bl_0_32 br_0_32 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c32
*+ bl_0_32 br_0_32 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c32
*+ bl_0_32 br_0_32 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c32
*+ bl_0_32 br_0_32 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c32
*+ bl_0_32 br_0_32 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c32
*+ bl_0_32 br_0_32 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c32
*+ bl_0_32 br_0_32 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c32
*+ bl_0_32 br_0_32 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c32
*+ bl_0_32 br_0_32 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c32
*+ bl_0_32 br_0_32 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c32
*+ bl_0_32 br_0_32 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c32
*+ bl_0_32 br_0_32 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c32
*+ bl_0_32 br_0_32 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c32
*+ bl_0_32 br_0_32 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c32
*+ bl_0_32 br_0_32 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c32
*+ bl_0_32 br_0_32 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c32
*+ bl_0_32 br_0_32 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c32
*+ bl_0_32 br_0_32 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c32
*+ bl_0_32 br_0_32 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c32
*+ bl_0_32 br_0_32 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c32
*+ bl_0_32 br_0_32 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c32
*+ bl_0_32 br_0_32 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c32
*+ bl_0_32 br_0_32 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c32
*+ bl_0_32 br_0_32 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c32
+ bl_0_32 br_0_32 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c33
*+ bl_0_33 br_0_33 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c33
*+ bl_0_33 br_0_33 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c33
*+ bl_0_33 br_0_33 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c33
*+ bl_0_33 br_0_33 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c33
*+ bl_0_33 br_0_33 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c33
*+ bl_0_33 br_0_33 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c33
*+ bl_0_33 br_0_33 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c33
*+ bl_0_33 br_0_33 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c33
*+ bl_0_33 br_0_33 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c33
*+ bl_0_33 br_0_33 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c33
*+ bl_0_33 br_0_33 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c33
*+ bl_0_33 br_0_33 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c33
*+ bl_0_33 br_0_33 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c33
*+ bl_0_33 br_0_33 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c33
*+ bl_0_33 br_0_33 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c33
*+ bl_0_33 br_0_33 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c33
*+ bl_0_33 br_0_33 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c33
*+ bl_0_33 br_0_33 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c33
*+ bl_0_33 br_0_33 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c33
*+ bl_0_33 br_0_33 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c33
*+ bl_0_33 br_0_33 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c33
*+ bl_0_33 br_0_33 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c33
*+ bl_0_33 br_0_33 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c33
*+ bl_0_33 br_0_33 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c33
*+ bl_0_33 br_0_33 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c33
*+ bl_0_33 br_0_33 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c33
*+ bl_0_33 br_0_33 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c33
*+ bl_0_33 br_0_33 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c33
*+ bl_0_33 br_0_33 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c33
*+ bl_0_33 br_0_33 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c33
+ bl_0_33 br_0_33 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c34
*+ bl_0_34 br_0_34 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c34
*+ bl_0_34 br_0_34 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c34
*+ bl_0_34 br_0_34 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c34
*+ bl_0_34 br_0_34 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c34
*+ bl_0_34 br_0_34 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c34
*+ bl_0_34 br_0_34 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c34
*+ bl_0_34 br_0_34 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c34
*+ bl_0_34 br_0_34 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c34
*+ bl_0_34 br_0_34 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c34
*+ bl_0_34 br_0_34 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c34
*+ bl_0_34 br_0_34 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c34
*+ bl_0_34 br_0_34 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c34
*+ bl_0_34 br_0_34 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c34
*+ bl_0_34 br_0_34 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c34
*+ bl_0_34 br_0_34 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c34
*+ bl_0_34 br_0_34 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c34
*+ bl_0_34 br_0_34 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c34
*+ bl_0_34 br_0_34 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c34
*+ bl_0_34 br_0_34 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c34
*+ bl_0_34 br_0_34 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c34
*+ bl_0_34 br_0_34 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c34
*+ bl_0_34 br_0_34 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c34
*+ bl_0_34 br_0_34 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c34
*+ bl_0_34 br_0_34 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c34
*+ bl_0_34 br_0_34 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c34
*+ bl_0_34 br_0_34 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c34
*+ bl_0_34 br_0_34 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c34
*+ bl_0_34 br_0_34 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c34
*+ bl_0_34 br_0_34 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c34
*+ bl_0_34 br_0_34 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c34
+ bl_0_34 br_0_34 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c35
*+ bl_0_35 br_0_35 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c35
*+ bl_0_35 br_0_35 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c35
*+ bl_0_35 br_0_35 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c35
*+ bl_0_35 br_0_35 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c35
*+ bl_0_35 br_0_35 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c35
*+ bl_0_35 br_0_35 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c35
*+ bl_0_35 br_0_35 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c35
*+ bl_0_35 br_0_35 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c35
*+ bl_0_35 br_0_35 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c35
*+ bl_0_35 br_0_35 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c35
*+ bl_0_35 br_0_35 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c35
*+ bl_0_35 br_0_35 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c35
*+ bl_0_35 br_0_35 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c35
*+ bl_0_35 br_0_35 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c35
*+ bl_0_35 br_0_35 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c35
*+ bl_0_35 br_0_35 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c35
*+ bl_0_35 br_0_35 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c35
*+ bl_0_35 br_0_35 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c35
*+ bl_0_35 br_0_35 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c35
*+ bl_0_35 br_0_35 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c35
*+ bl_0_35 br_0_35 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c35
*+ bl_0_35 br_0_35 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c35
*+ bl_0_35 br_0_35 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c35
*+ bl_0_35 br_0_35 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c35
*+ bl_0_35 br_0_35 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c35
*+ bl_0_35 br_0_35 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c35
*+ bl_0_35 br_0_35 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c35
*+ bl_0_35 br_0_35 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c35
*+ bl_0_35 br_0_35 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c35
*+ bl_0_35 br_0_35 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c35
+ bl_0_35 br_0_35 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c36
*+ bl_0_36 br_0_36 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c36
*+ bl_0_36 br_0_36 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c36
*+ bl_0_36 br_0_36 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c36
*+ bl_0_36 br_0_36 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c36
*+ bl_0_36 br_0_36 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c36
*+ bl_0_36 br_0_36 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c36
*+ bl_0_36 br_0_36 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c36
*+ bl_0_36 br_0_36 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c36
*+ bl_0_36 br_0_36 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c36
*+ bl_0_36 br_0_36 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c36
*+ bl_0_36 br_0_36 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c36
*+ bl_0_36 br_0_36 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c36
*+ bl_0_36 br_0_36 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c36
*+ bl_0_36 br_0_36 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c36
*+ bl_0_36 br_0_36 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c36
*+ bl_0_36 br_0_36 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c36
*+ bl_0_36 br_0_36 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c36
*+ bl_0_36 br_0_36 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c36
*+ bl_0_36 br_0_36 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c36
*+ bl_0_36 br_0_36 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c36
*+ bl_0_36 br_0_36 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c36
*+ bl_0_36 br_0_36 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c36
*+ bl_0_36 br_0_36 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c36
*+ bl_0_36 br_0_36 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c36
*+ bl_0_36 br_0_36 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c36
*+ bl_0_36 br_0_36 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c36
*+ bl_0_36 br_0_36 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c36
*+ bl_0_36 br_0_36 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c36
*+ bl_0_36 br_0_36 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c36
*+ bl_0_36 br_0_36 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c36
+ bl_0_36 br_0_36 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c37
*+ bl_0_37 br_0_37 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c37
*+ bl_0_37 br_0_37 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c37
*+ bl_0_37 br_0_37 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c37
*+ bl_0_37 br_0_37 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c37
*+ bl_0_37 br_0_37 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c37
*+ bl_0_37 br_0_37 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c37
*+ bl_0_37 br_0_37 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c37
*+ bl_0_37 br_0_37 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c37
*+ bl_0_37 br_0_37 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c37
*+ bl_0_37 br_0_37 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c37
*+ bl_0_37 br_0_37 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c37
*+ bl_0_37 br_0_37 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c37
*+ bl_0_37 br_0_37 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c37
*+ bl_0_37 br_0_37 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c37
*+ bl_0_37 br_0_37 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c37
*+ bl_0_37 br_0_37 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c37
*+ bl_0_37 br_0_37 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c37
*+ bl_0_37 br_0_37 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c37
*+ bl_0_37 br_0_37 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c37
*+ bl_0_37 br_0_37 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c37
*+ bl_0_37 br_0_37 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c37
*+ bl_0_37 br_0_37 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c37
*+ bl_0_37 br_0_37 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c37
*+ bl_0_37 br_0_37 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c37
*+ bl_0_37 br_0_37 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c37
*+ bl_0_37 br_0_37 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c37
*+ bl_0_37 br_0_37 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c37
*+ bl_0_37 br_0_37 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c37
*+ bl_0_37 br_0_37 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c37
*+ bl_0_37 br_0_37 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c37
+ bl_0_37 br_0_37 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c38
*+ bl_0_38 br_0_38 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c38
*+ bl_0_38 br_0_38 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c38
*+ bl_0_38 br_0_38 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c38
*+ bl_0_38 br_0_38 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c38
*+ bl_0_38 br_0_38 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c38
*+ bl_0_38 br_0_38 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c38
*+ bl_0_38 br_0_38 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c38
*+ bl_0_38 br_0_38 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c38
*+ bl_0_38 br_0_38 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c38
*+ bl_0_38 br_0_38 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c38
*+ bl_0_38 br_0_38 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c38
*+ bl_0_38 br_0_38 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c38
*+ bl_0_38 br_0_38 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c38
*+ bl_0_38 br_0_38 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c38
*+ bl_0_38 br_0_38 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c38
*+ bl_0_38 br_0_38 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c38
*+ bl_0_38 br_0_38 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c38
*+ bl_0_38 br_0_38 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c38
*+ bl_0_38 br_0_38 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c38
*+ bl_0_38 br_0_38 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c38
*+ bl_0_38 br_0_38 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c38
*+ bl_0_38 br_0_38 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c38
*+ bl_0_38 br_0_38 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c38
*+ bl_0_38 br_0_38 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c38
*+ bl_0_38 br_0_38 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c38
*+ bl_0_38 br_0_38 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c38
*+ bl_0_38 br_0_38 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c38
*+ bl_0_38 br_0_38 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c38
*+ bl_0_38 br_0_38 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c38
*+ bl_0_38 br_0_38 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c38
+ bl_0_38 br_0_38 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c39
*+ bl_0_39 br_0_39 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c39
*+ bl_0_39 br_0_39 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c39
*+ bl_0_39 br_0_39 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c39
*+ bl_0_39 br_0_39 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c39
*+ bl_0_39 br_0_39 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c39
*+ bl_0_39 br_0_39 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c39
*+ bl_0_39 br_0_39 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c39
*+ bl_0_39 br_0_39 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c39
*+ bl_0_39 br_0_39 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c39
*+ bl_0_39 br_0_39 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c39
*+ bl_0_39 br_0_39 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c39
*+ bl_0_39 br_0_39 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c39
*+ bl_0_39 br_0_39 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c39
*+ bl_0_39 br_0_39 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c39
*+ bl_0_39 br_0_39 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c39
*+ bl_0_39 br_0_39 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c39
*+ bl_0_39 br_0_39 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c39
*+ bl_0_39 br_0_39 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c39
*+ bl_0_39 br_0_39 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c39
*+ bl_0_39 br_0_39 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c39
*+ bl_0_39 br_0_39 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c39
*+ bl_0_39 br_0_39 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c39
*+ bl_0_39 br_0_39 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c39
*+ bl_0_39 br_0_39 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c39
*+ bl_0_39 br_0_39 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c39
*+ bl_0_39 br_0_39 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c39
*+ bl_0_39 br_0_39 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c39
*+ bl_0_39 br_0_39 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c39
*+ bl_0_39 br_0_39 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c39
*+ bl_0_39 br_0_39 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c39
+ bl_0_39 br_0_39 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c40
*+ bl_0_40 br_0_40 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c40
*+ bl_0_40 br_0_40 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c40
*+ bl_0_40 br_0_40 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c40
*+ bl_0_40 br_0_40 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c40
*+ bl_0_40 br_0_40 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c40
*+ bl_0_40 br_0_40 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c40
*+ bl_0_40 br_0_40 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c40
*+ bl_0_40 br_0_40 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c40
*+ bl_0_40 br_0_40 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c40
*+ bl_0_40 br_0_40 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c40
*+ bl_0_40 br_0_40 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c40
*+ bl_0_40 br_0_40 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c40
*+ bl_0_40 br_0_40 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c40
*+ bl_0_40 br_0_40 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c40
*+ bl_0_40 br_0_40 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c40
*+ bl_0_40 br_0_40 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c40
*+ bl_0_40 br_0_40 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c40
*+ bl_0_40 br_0_40 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c40
*+ bl_0_40 br_0_40 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c40
*+ bl_0_40 br_0_40 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c40
*+ bl_0_40 br_0_40 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c40
*+ bl_0_40 br_0_40 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c40
*+ bl_0_40 br_0_40 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c40
*+ bl_0_40 br_0_40 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c40
*+ bl_0_40 br_0_40 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c40
*+ bl_0_40 br_0_40 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c40
*+ bl_0_40 br_0_40 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c40
*+ bl_0_40 br_0_40 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c40
*+ bl_0_40 br_0_40 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c40
*+ bl_0_40 br_0_40 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c40
+ bl_0_40 br_0_40 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c41
*+ bl_0_41 br_0_41 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c41
*+ bl_0_41 br_0_41 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c41
*+ bl_0_41 br_0_41 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c41
*+ bl_0_41 br_0_41 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c41
*+ bl_0_41 br_0_41 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c41
*+ bl_0_41 br_0_41 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c41
*+ bl_0_41 br_0_41 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c41
*+ bl_0_41 br_0_41 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c41
*+ bl_0_41 br_0_41 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c41
*+ bl_0_41 br_0_41 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c41
*+ bl_0_41 br_0_41 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c41
*+ bl_0_41 br_0_41 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c41
*+ bl_0_41 br_0_41 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c41
*+ bl_0_41 br_0_41 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c41
*+ bl_0_41 br_0_41 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c41
*+ bl_0_41 br_0_41 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c41
*+ bl_0_41 br_0_41 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c41
*+ bl_0_41 br_0_41 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c41
*+ bl_0_41 br_0_41 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c41
*+ bl_0_41 br_0_41 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c41
*+ bl_0_41 br_0_41 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c41
*+ bl_0_41 br_0_41 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c41
*+ bl_0_41 br_0_41 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c41
*+ bl_0_41 br_0_41 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c41
*+ bl_0_41 br_0_41 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c41
*+ bl_0_41 br_0_41 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c41
*+ bl_0_41 br_0_41 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c41
*+ bl_0_41 br_0_41 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c41
*+ bl_0_41 br_0_41 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c41
*+ bl_0_41 br_0_41 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c41
+ bl_0_41 br_0_41 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c42
*+ bl_0_42 br_0_42 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c42
*+ bl_0_42 br_0_42 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c42
*+ bl_0_42 br_0_42 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c42
*+ bl_0_42 br_0_42 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c42
*+ bl_0_42 br_0_42 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c42
*+ bl_0_42 br_0_42 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c42
*+ bl_0_42 br_0_42 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c42
*+ bl_0_42 br_0_42 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c42
*+ bl_0_42 br_0_42 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c42
*+ bl_0_42 br_0_42 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c42
*+ bl_0_42 br_0_42 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c42
*+ bl_0_42 br_0_42 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c42
*+ bl_0_42 br_0_42 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c42
*+ bl_0_42 br_0_42 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c42
*+ bl_0_42 br_0_42 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c42
*+ bl_0_42 br_0_42 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c42
*+ bl_0_42 br_0_42 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c42
*+ bl_0_42 br_0_42 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c42
*+ bl_0_42 br_0_42 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c42
*+ bl_0_42 br_0_42 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c42
*+ bl_0_42 br_0_42 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c42
*+ bl_0_42 br_0_42 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c42
*+ bl_0_42 br_0_42 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c42
*+ bl_0_42 br_0_42 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c42
*+ bl_0_42 br_0_42 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c42
*+ bl_0_42 br_0_42 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c42
*+ bl_0_42 br_0_42 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c42
*+ bl_0_42 br_0_42 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c42
*+ bl_0_42 br_0_42 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c42
*+ bl_0_42 br_0_42 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c42
+ bl_0_42 br_0_42 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c43
*+ bl_0_43 br_0_43 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c43
*+ bl_0_43 br_0_43 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c43
*+ bl_0_43 br_0_43 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c43
*+ bl_0_43 br_0_43 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c43
*+ bl_0_43 br_0_43 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c43
*+ bl_0_43 br_0_43 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c43
*+ bl_0_43 br_0_43 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c43
*+ bl_0_43 br_0_43 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c43
*+ bl_0_43 br_0_43 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c43
*+ bl_0_43 br_0_43 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c43
*+ bl_0_43 br_0_43 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c43
*+ bl_0_43 br_0_43 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c43
*+ bl_0_43 br_0_43 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c43
*+ bl_0_43 br_0_43 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c43
*+ bl_0_43 br_0_43 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c43
*+ bl_0_43 br_0_43 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c43
*+ bl_0_43 br_0_43 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c43
*+ bl_0_43 br_0_43 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c43
*+ bl_0_43 br_0_43 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c43
*+ bl_0_43 br_0_43 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c43
*+ bl_0_43 br_0_43 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c43
*+ bl_0_43 br_0_43 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c43
*+ bl_0_43 br_0_43 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c43
*+ bl_0_43 br_0_43 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c43
*+ bl_0_43 br_0_43 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c43
*+ bl_0_43 br_0_43 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c43
*+ bl_0_43 br_0_43 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c43
*+ bl_0_43 br_0_43 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c43
*+ bl_0_43 br_0_43 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c43
*+ bl_0_43 br_0_43 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c43
+ bl_0_43 br_0_43 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c44
*+ bl_0_44 br_0_44 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c44
*+ bl_0_44 br_0_44 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c44
*+ bl_0_44 br_0_44 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c44
*+ bl_0_44 br_0_44 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c44
*+ bl_0_44 br_0_44 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c44
*+ bl_0_44 br_0_44 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c44
*+ bl_0_44 br_0_44 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c44
*+ bl_0_44 br_0_44 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c44
*+ bl_0_44 br_0_44 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c44
*+ bl_0_44 br_0_44 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c44
*+ bl_0_44 br_0_44 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c44
*+ bl_0_44 br_0_44 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c44
*+ bl_0_44 br_0_44 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c44
*+ bl_0_44 br_0_44 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c44
*+ bl_0_44 br_0_44 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c44
*+ bl_0_44 br_0_44 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c44
*+ bl_0_44 br_0_44 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c44
*+ bl_0_44 br_0_44 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c44
*+ bl_0_44 br_0_44 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c44
*+ bl_0_44 br_0_44 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c44
*+ bl_0_44 br_0_44 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c44
*+ bl_0_44 br_0_44 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c44
*+ bl_0_44 br_0_44 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c44
*+ bl_0_44 br_0_44 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c44
*+ bl_0_44 br_0_44 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c44
*+ bl_0_44 br_0_44 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c44
*+ bl_0_44 br_0_44 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c44
*+ bl_0_44 br_0_44 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c44
*+ bl_0_44 br_0_44 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c44
*+ bl_0_44 br_0_44 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c44
+ bl_0_44 br_0_44 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c45
*+ bl_0_45 br_0_45 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c45
*+ bl_0_45 br_0_45 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c45
*+ bl_0_45 br_0_45 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c45
*+ bl_0_45 br_0_45 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c45
*+ bl_0_45 br_0_45 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c45
*+ bl_0_45 br_0_45 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c45
*+ bl_0_45 br_0_45 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c45
*+ bl_0_45 br_0_45 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c45
*+ bl_0_45 br_0_45 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c45
*+ bl_0_45 br_0_45 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c45
*+ bl_0_45 br_0_45 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c45
*+ bl_0_45 br_0_45 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c45
*+ bl_0_45 br_0_45 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c45
*+ bl_0_45 br_0_45 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c45
*+ bl_0_45 br_0_45 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c45
*+ bl_0_45 br_0_45 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c45
*+ bl_0_45 br_0_45 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c45
*+ bl_0_45 br_0_45 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c45
*+ bl_0_45 br_0_45 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c45
*+ bl_0_45 br_0_45 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c45
*+ bl_0_45 br_0_45 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c45
*+ bl_0_45 br_0_45 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c45
*+ bl_0_45 br_0_45 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c45
*+ bl_0_45 br_0_45 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c45
*+ bl_0_45 br_0_45 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c45
*+ bl_0_45 br_0_45 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c45
*+ bl_0_45 br_0_45 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c45
*+ bl_0_45 br_0_45 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c45
*+ bl_0_45 br_0_45 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c45
*+ bl_0_45 br_0_45 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c45
+ bl_0_45 br_0_45 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c46
*+ bl_0_46 br_0_46 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c46
*+ bl_0_46 br_0_46 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c46
*+ bl_0_46 br_0_46 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c46
*+ bl_0_46 br_0_46 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c46
*+ bl_0_46 br_0_46 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c46
*+ bl_0_46 br_0_46 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c46
*+ bl_0_46 br_0_46 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c46
*+ bl_0_46 br_0_46 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c46
*+ bl_0_46 br_0_46 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c46
*+ bl_0_46 br_0_46 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c46
*+ bl_0_46 br_0_46 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c46
*+ bl_0_46 br_0_46 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c46
*+ bl_0_46 br_0_46 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c46
*+ bl_0_46 br_0_46 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c46
*+ bl_0_46 br_0_46 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c46
*+ bl_0_46 br_0_46 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c46
*+ bl_0_46 br_0_46 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c46
*+ bl_0_46 br_0_46 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c46
*+ bl_0_46 br_0_46 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c46
*+ bl_0_46 br_0_46 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c46
*+ bl_0_46 br_0_46 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c46
*+ bl_0_46 br_0_46 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c46
*+ bl_0_46 br_0_46 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c46
*+ bl_0_46 br_0_46 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c46
*+ bl_0_46 br_0_46 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c46
*+ bl_0_46 br_0_46 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c46
*+ bl_0_46 br_0_46 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c46
*+ bl_0_46 br_0_46 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c46
*+ bl_0_46 br_0_46 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c46
*+ bl_0_46 br_0_46 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c46
+ bl_0_46 br_0_46 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c47
*+ bl_0_47 br_0_47 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c47
*+ bl_0_47 br_0_47 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c47
*+ bl_0_47 br_0_47 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c47
*+ bl_0_47 br_0_47 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c47
*+ bl_0_47 br_0_47 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c47
*+ bl_0_47 br_0_47 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c47
*+ bl_0_47 br_0_47 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c47
*+ bl_0_47 br_0_47 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c47
*+ bl_0_47 br_0_47 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c47
*+ bl_0_47 br_0_47 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c47
*+ bl_0_47 br_0_47 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c47
*+ bl_0_47 br_0_47 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c47
*+ bl_0_47 br_0_47 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c47
*+ bl_0_47 br_0_47 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c47
*+ bl_0_47 br_0_47 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c47
*+ bl_0_47 br_0_47 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c47
*+ bl_0_47 br_0_47 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c47
*+ bl_0_47 br_0_47 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c47
*+ bl_0_47 br_0_47 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c47
*+ bl_0_47 br_0_47 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c47
*+ bl_0_47 br_0_47 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c47
*+ bl_0_47 br_0_47 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c47
*+ bl_0_47 br_0_47 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c47
*+ bl_0_47 br_0_47 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c47
*+ bl_0_47 br_0_47 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c47
*+ bl_0_47 br_0_47 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c47
*+ bl_0_47 br_0_47 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c47
*+ bl_0_47 br_0_47 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c47
*+ bl_0_47 br_0_47 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c47
*+ bl_0_47 br_0_47 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c47
+ bl_0_47 br_0_47 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c48
*+ bl_0_48 br_0_48 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c48
*+ bl_0_48 br_0_48 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c48
*+ bl_0_48 br_0_48 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c48
*+ bl_0_48 br_0_48 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c48
*+ bl_0_48 br_0_48 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c48
*+ bl_0_48 br_0_48 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c48
*+ bl_0_48 br_0_48 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c48
*+ bl_0_48 br_0_48 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c48
*+ bl_0_48 br_0_48 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c48
*+ bl_0_48 br_0_48 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c48
*+ bl_0_48 br_0_48 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c48
*+ bl_0_48 br_0_48 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c48
*+ bl_0_48 br_0_48 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c48
*+ bl_0_48 br_0_48 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c48
*+ bl_0_48 br_0_48 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c48
*+ bl_0_48 br_0_48 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c48
*+ bl_0_48 br_0_48 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c48
*+ bl_0_48 br_0_48 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c48
*+ bl_0_48 br_0_48 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c48
*+ bl_0_48 br_0_48 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c48
*+ bl_0_48 br_0_48 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c48
*+ bl_0_48 br_0_48 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c48
*+ bl_0_48 br_0_48 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c48
*+ bl_0_48 br_0_48 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c48
*+ bl_0_48 br_0_48 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c48
*+ bl_0_48 br_0_48 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c48
*+ bl_0_48 br_0_48 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c48
*+ bl_0_48 br_0_48 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c48
*+ bl_0_48 br_0_48 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c48
*+ bl_0_48 br_0_48 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c48
+ bl_0_48 br_0_48 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c49
*+ bl_0_49 br_0_49 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c49
*+ bl_0_49 br_0_49 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c49
*+ bl_0_49 br_0_49 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c49
*+ bl_0_49 br_0_49 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c49
*+ bl_0_49 br_0_49 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c49
*+ bl_0_49 br_0_49 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c49
*+ bl_0_49 br_0_49 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c49
*+ bl_0_49 br_0_49 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c49
*+ bl_0_49 br_0_49 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c49
*+ bl_0_49 br_0_49 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c49
*+ bl_0_49 br_0_49 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c49
*+ bl_0_49 br_0_49 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c49
*+ bl_0_49 br_0_49 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c49
*+ bl_0_49 br_0_49 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c49
*+ bl_0_49 br_0_49 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c49
*+ bl_0_49 br_0_49 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c49
*+ bl_0_49 br_0_49 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c49
*+ bl_0_49 br_0_49 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c49
*+ bl_0_49 br_0_49 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c49
*+ bl_0_49 br_0_49 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c49
*+ bl_0_49 br_0_49 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c49
*+ bl_0_49 br_0_49 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c49
*+ bl_0_49 br_0_49 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c49
*+ bl_0_49 br_0_49 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c49
*+ bl_0_49 br_0_49 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c49
*+ bl_0_49 br_0_49 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c49
*+ bl_0_49 br_0_49 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c49
*+ bl_0_49 br_0_49 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c49
*+ bl_0_49 br_0_49 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c49
*+ bl_0_49 br_0_49 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c49
+ bl_0_49 br_0_49 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c50
*+ bl_0_50 br_0_50 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c50
*+ bl_0_50 br_0_50 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c50
*+ bl_0_50 br_0_50 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c50
*+ bl_0_50 br_0_50 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c50
*+ bl_0_50 br_0_50 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c50
*+ bl_0_50 br_0_50 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c50
*+ bl_0_50 br_0_50 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c50
*+ bl_0_50 br_0_50 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c50
*+ bl_0_50 br_0_50 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c50
*+ bl_0_50 br_0_50 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c50
*+ bl_0_50 br_0_50 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c50
*+ bl_0_50 br_0_50 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c50
*+ bl_0_50 br_0_50 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c50
*+ bl_0_50 br_0_50 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c50
*+ bl_0_50 br_0_50 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c50
*+ bl_0_50 br_0_50 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c50
*+ bl_0_50 br_0_50 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c50
*+ bl_0_50 br_0_50 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c50
*+ bl_0_50 br_0_50 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c50
*+ bl_0_50 br_0_50 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c50
*+ bl_0_50 br_0_50 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c50
*+ bl_0_50 br_0_50 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c50
*+ bl_0_50 br_0_50 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c50
*+ bl_0_50 br_0_50 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c50
*+ bl_0_50 br_0_50 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c50
*+ bl_0_50 br_0_50 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c50
*+ bl_0_50 br_0_50 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c50
*+ bl_0_50 br_0_50 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c50
*+ bl_0_50 br_0_50 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c50
*+ bl_0_50 br_0_50 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c50
+ bl_0_50 br_0_50 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c51
*+ bl_0_51 br_0_51 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c51
*+ bl_0_51 br_0_51 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c51
*+ bl_0_51 br_0_51 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c51
*+ bl_0_51 br_0_51 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c51
*+ bl_0_51 br_0_51 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c51
*+ bl_0_51 br_0_51 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c51
*+ bl_0_51 br_0_51 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c51
*+ bl_0_51 br_0_51 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c51
*+ bl_0_51 br_0_51 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c51
*+ bl_0_51 br_0_51 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c51
*+ bl_0_51 br_0_51 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c51
*+ bl_0_51 br_0_51 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c51
*+ bl_0_51 br_0_51 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c51
*+ bl_0_51 br_0_51 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c51
*+ bl_0_51 br_0_51 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c51
*+ bl_0_51 br_0_51 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c51
*+ bl_0_51 br_0_51 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c51
*+ bl_0_51 br_0_51 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c51
*+ bl_0_51 br_0_51 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c51
*+ bl_0_51 br_0_51 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c51
*+ bl_0_51 br_0_51 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c51
*+ bl_0_51 br_0_51 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c51
*+ bl_0_51 br_0_51 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c51
*+ bl_0_51 br_0_51 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c51
*+ bl_0_51 br_0_51 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c51
*+ bl_0_51 br_0_51 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c51
*+ bl_0_51 br_0_51 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c51
*+ bl_0_51 br_0_51 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c51
*+ bl_0_51 br_0_51 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c51
*+ bl_0_51 br_0_51 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c51
+ bl_0_51 br_0_51 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c52
*+ bl_0_52 br_0_52 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c52
*+ bl_0_52 br_0_52 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c52
*+ bl_0_52 br_0_52 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c52
*+ bl_0_52 br_0_52 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c52
*+ bl_0_52 br_0_52 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c52
*+ bl_0_52 br_0_52 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c52
*+ bl_0_52 br_0_52 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c52
*+ bl_0_52 br_0_52 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c52
*+ bl_0_52 br_0_52 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c52
*+ bl_0_52 br_0_52 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c52
*+ bl_0_52 br_0_52 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c52
*+ bl_0_52 br_0_52 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c52
*+ bl_0_52 br_0_52 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c52
*+ bl_0_52 br_0_52 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c52
*+ bl_0_52 br_0_52 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c52
*+ bl_0_52 br_0_52 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c52
*+ bl_0_52 br_0_52 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c52
*+ bl_0_52 br_0_52 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c52
*+ bl_0_52 br_0_52 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c52
*+ bl_0_52 br_0_52 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c52
*+ bl_0_52 br_0_52 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c52
*+ bl_0_52 br_0_52 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c52
*+ bl_0_52 br_0_52 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c52
*+ bl_0_52 br_0_52 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c52
*+ bl_0_52 br_0_52 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c52
*+ bl_0_52 br_0_52 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c52
*+ bl_0_52 br_0_52 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c52
*+ bl_0_52 br_0_52 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c52
*+ bl_0_52 br_0_52 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c52
*+ bl_0_52 br_0_52 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c52
+ bl_0_52 br_0_52 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c53
*+ bl_0_53 br_0_53 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c53
*+ bl_0_53 br_0_53 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c53
*+ bl_0_53 br_0_53 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c53
*+ bl_0_53 br_0_53 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c53
*+ bl_0_53 br_0_53 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c53
*+ bl_0_53 br_0_53 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c53
*+ bl_0_53 br_0_53 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c53
*+ bl_0_53 br_0_53 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c53
*+ bl_0_53 br_0_53 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c53
*+ bl_0_53 br_0_53 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c53
*+ bl_0_53 br_0_53 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c53
*+ bl_0_53 br_0_53 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c53
*+ bl_0_53 br_0_53 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c53
*+ bl_0_53 br_0_53 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c53
*+ bl_0_53 br_0_53 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c53
*+ bl_0_53 br_0_53 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c53
*+ bl_0_53 br_0_53 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c53
*+ bl_0_53 br_0_53 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c53
*+ bl_0_53 br_0_53 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c53
*+ bl_0_53 br_0_53 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c53
*+ bl_0_53 br_0_53 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c53
*+ bl_0_53 br_0_53 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c53
*+ bl_0_53 br_0_53 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c53
*+ bl_0_53 br_0_53 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c53
*+ bl_0_53 br_0_53 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c53
*+ bl_0_53 br_0_53 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c53
*+ bl_0_53 br_0_53 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c53
*+ bl_0_53 br_0_53 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c53
*+ bl_0_53 br_0_53 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c53
*+ bl_0_53 br_0_53 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c53
+ bl_0_53 br_0_53 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c54
*+ bl_0_54 br_0_54 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c54
*+ bl_0_54 br_0_54 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c54
*+ bl_0_54 br_0_54 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c54
*+ bl_0_54 br_0_54 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c54
*+ bl_0_54 br_0_54 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c54
*+ bl_0_54 br_0_54 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c54
*+ bl_0_54 br_0_54 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c54
*+ bl_0_54 br_0_54 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c54
*+ bl_0_54 br_0_54 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c54
*+ bl_0_54 br_0_54 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c54
*+ bl_0_54 br_0_54 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c54
*+ bl_0_54 br_0_54 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c54
*+ bl_0_54 br_0_54 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c54
*+ bl_0_54 br_0_54 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c54
*+ bl_0_54 br_0_54 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c54
*+ bl_0_54 br_0_54 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c54
*+ bl_0_54 br_0_54 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c54
*+ bl_0_54 br_0_54 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c54
*+ bl_0_54 br_0_54 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c54
*+ bl_0_54 br_0_54 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c54
*+ bl_0_54 br_0_54 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c54
*+ bl_0_54 br_0_54 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c54
*+ bl_0_54 br_0_54 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c54
*+ bl_0_54 br_0_54 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c54
*+ bl_0_54 br_0_54 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c54
*+ bl_0_54 br_0_54 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c54
*+ bl_0_54 br_0_54 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c54
*+ bl_0_54 br_0_54 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c54
*+ bl_0_54 br_0_54 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c54
*+ bl_0_54 br_0_54 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c54
+ bl_0_54 br_0_54 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c55
*+ bl_0_55 br_0_55 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c55
*+ bl_0_55 br_0_55 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c55
*+ bl_0_55 br_0_55 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c55
*+ bl_0_55 br_0_55 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c55
*+ bl_0_55 br_0_55 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c55
*+ bl_0_55 br_0_55 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c55
*+ bl_0_55 br_0_55 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c55
*+ bl_0_55 br_0_55 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c55
*+ bl_0_55 br_0_55 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c55
*+ bl_0_55 br_0_55 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c55
*+ bl_0_55 br_0_55 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c55
*+ bl_0_55 br_0_55 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c55
*+ bl_0_55 br_0_55 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c55
*+ bl_0_55 br_0_55 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c55
*+ bl_0_55 br_0_55 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c55
*+ bl_0_55 br_0_55 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c55
*+ bl_0_55 br_0_55 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c55
*+ bl_0_55 br_0_55 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c55
*+ bl_0_55 br_0_55 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c55
*+ bl_0_55 br_0_55 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c55
*+ bl_0_55 br_0_55 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c55
*+ bl_0_55 br_0_55 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c55
*+ bl_0_55 br_0_55 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c55
*+ bl_0_55 br_0_55 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c55
*+ bl_0_55 br_0_55 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c55
*+ bl_0_55 br_0_55 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c55
*+ bl_0_55 br_0_55 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c55
*+ bl_0_55 br_0_55 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c55
*+ bl_0_55 br_0_55 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c55
*+ bl_0_55 br_0_55 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c55
+ bl_0_55 br_0_55 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c56
*+ bl_0_56 br_0_56 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c56
*+ bl_0_56 br_0_56 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c56
*+ bl_0_56 br_0_56 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c56
*+ bl_0_56 br_0_56 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c56
*+ bl_0_56 br_0_56 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c56
*+ bl_0_56 br_0_56 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c56
*+ bl_0_56 br_0_56 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c56
*+ bl_0_56 br_0_56 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c56
*+ bl_0_56 br_0_56 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c56
*+ bl_0_56 br_0_56 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c56
*+ bl_0_56 br_0_56 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c56
*+ bl_0_56 br_0_56 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c56
*+ bl_0_56 br_0_56 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c56
*+ bl_0_56 br_0_56 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c56
*+ bl_0_56 br_0_56 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c56
*+ bl_0_56 br_0_56 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c56
*+ bl_0_56 br_0_56 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c56
*+ bl_0_56 br_0_56 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c56
*+ bl_0_56 br_0_56 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c56
*+ bl_0_56 br_0_56 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c56
*+ bl_0_56 br_0_56 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c56
*+ bl_0_56 br_0_56 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c56
*+ bl_0_56 br_0_56 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c56
*+ bl_0_56 br_0_56 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c56
*+ bl_0_56 br_0_56 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c56
*+ bl_0_56 br_0_56 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c56
*+ bl_0_56 br_0_56 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c56
*+ bl_0_56 br_0_56 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c56
*+ bl_0_56 br_0_56 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c56
*+ bl_0_56 br_0_56 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c56
+ bl_0_56 br_0_56 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c57
*+ bl_0_57 br_0_57 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c57
*+ bl_0_57 br_0_57 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c57
*+ bl_0_57 br_0_57 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c57
*+ bl_0_57 br_0_57 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c57
*+ bl_0_57 br_0_57 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c57
*+ bl_0_57 br_0_57 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c57
*+ bl_0_57 br_0_57 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c57
*+ bl_0_57 br_0_57 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c57
*+ bl_0_57 br_0_57 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c57
*+ bl_0_57 br_0_57 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c57
*+ bl_0_57 br_0_57 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c57
*+ bl_0_57 br_0_57 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c57
*+ bl_0_57 br_0_57 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c57
*+ bl_0_57 br_0_57 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c57
*+ bl_0_57 br_0_57 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c57
*+ bl_0_57 br_0_57 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c57
*+ bl_0_57 br_0_57 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c57
*+ bl_0_57 br_0_57 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c57
*+ bl_0_57 br_0_57 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c57
*+ bl_0_57 br_0_57 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c57
*+ bl_0_57 br_0_57 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c57
*+ bl_0_57 br_0_57 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c57
*+ bl_0_57 br_0_57 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c57
*+ bl_0_57 br_0_57 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c57
*+ bl_0_57 br_0_57 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c57
*+ bl_0_57 br_0_57 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c57
*+ bl_0_57 br_0_57 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c57
*+ bl_0_57 br_0_57 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c57
*+ bl_0_57 br_0_57 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c57
*+ bl_0_57 br_0_57 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c57
+ bl_0_57 br_0_57 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c58
*+ bl_0_58 br_0_58 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c58
*+ bl_0_58 br_0_58 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c58
*+ bl_0_58 br_0_58 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c58
*+ bl_0_58 br_0_58 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c58
*+ bl_0_58 br_0_58 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c58
*+ bl_0_58 br_0_58 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c58
*+ bl_0_58 br_0_58 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c58
*+ bl_0_58 br_0_58 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c58
*+ bl_0_58 br_0_58 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c58
*+ bl_0_58 br_0_58 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c58
*+ bl_0_58 br_0_58 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c58
*+ bl_0_58 br_0_58 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c58
*+ bl_0_58 br_0_58 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c58
*+ bl_0_58 br_0_58 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c58
*+ bl_0_58 br_0_58 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c58
*+ bl_0_58 br_0_58 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c58
*+ bl_0_58 br_0_58 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c58
*+ bl_0_58 br_0_58 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c58
*+ bl_0_58 br_0_58 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c58
*+ bl_0_58 br_0_58 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c58
*+ bl_0_58 br_0_58 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c58
*+ bl_0_58 br_0_58 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c58
*+ bl_0_58 br_0_58 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c58
*+ bl_0_58 br_0_58 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c58
*+ bl_0_58 br_0_58 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c58
*+ bl_0_58 br_0_58 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c58
*+ bl_0_58 br_0_58 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c58
*+ bl_0_58 br_0_58 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c58
*+ bl_0_58 br_0_58 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c58
*+ bl_0_58 br_0_58 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c58
+ bl_0_58 br_0_58 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c59
*+ bl_0_59 br_0_59 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c59
*+ bl_0_59 br_0_59 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c59
*+ bl_0_59 br_0_59 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c59
*+ bl_0_59 br_0_59 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c59
*+ bl_0_59 br_0_59 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c59
*+ bl_0_59 br_0_59 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c59
*+ bl_0_59 br_0_59 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c59
*+ bl_0_59 br_0_59 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c59
*+ bl_0_59 br_0_59 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c59
*+ bl_0_59 br_0_59 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c59
*+ bl_0_59 br_0_59 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c59
*+ bl_0_59 br_0_59 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c59
*+ bl_0_59 br_0_59 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c59
*+ bl_0_59 br_0_59 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c59
*+ bl_0_59 br_0_59 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c59
*+ bl_0_59 br_0_59 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c59
*+ bl_0_59 br_0_59 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c59
*+ bl_0_59 br_0_59 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c59
*+ bl_0_59 br_0_59 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c59
*+ bl_0_59 br_0_59 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c59
*+ bl_0_59 br_0_59 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c59
*+ bl_0_59 br_0_59 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c59
*+ bl_0_59 br_0_59 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c59
*+ bl_0_59 br_0_59 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c59
*+ bl_0_59 br_0_59 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c59
*+ bl_0_59 br_0_59 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c59
*+ bl_0_59 br_0_59 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c59
*+ bl_0_59 br_0_59 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c59
*+ bl_0_59 br_0_59 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c59
*+ bl_0_59 br_0_59 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c59
+ bl_0_59 br_0_59 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c60
*+ bl_0_60 br_0_60 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c60
*+ bl_0_60 br_0_60 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c60
*+ bl_0_60 br_0_60 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c60
*+ bl_0_60 br_0_60 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c60
*+ bl_0_60 br_0_60 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c60
*+ bl_0_60 br_0_60 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c60
*+ bl_0_60 br_0_60 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c60
*+ bl_0_60 br_0_60 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c60
*+ bl_0_60 br_0_60 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c60
*+ bl_0_60 br_0_60 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c60
*+ bl_0_60 br_0_60 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c60
*+ bl_0_60 br_0_60 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c60
*+ bl_0_60 br_0_60 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c60
*+ bl_0_60 br_0_60 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c60
*+ bl_0_60 br_0_60 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c60
*+ bl_0_60 br_0_60 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c60
*+ bl_0_60 br_0_60 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c60
*+ bl_0_60 br_0_60 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c60
*+ bl_0_60 br_0_60 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c60
*+ bl_0_60 br_0_60 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c60
*+ bl_0_60 br_0_60 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c60
*+ bl_0_60 br_0_60 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c60
*+ bl_0_60 br_0_60 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c60
*+ bl_0_60 br_0_60 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c60
*+ bl_0_60 br_0_60 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c60
*+ bl_0_60 br_0_60 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c60
*+ bl_0_60 br_0_60 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c60
*+ bl_0_60 br_0_60 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c60
*+ bl_0_60 br_0_60 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c60
*+ bl_0_60 br_0_60 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c60
+ bl_0_60 br_0_60 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c61
*+ bl_0_61 br_0_61 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c61
*+ bl_0_61 br_0_61 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c61
*+ bl_0_61 br_0_61 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c61
*+ bl_0_61 br_0_61 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c61
*+ bl_0_61 br_0_61 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c61
*+ bl_0_61 br_0_61 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c61
*+ bl_0_61 br_0_61 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c61
*+ bl_0_61 br_0_61 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c61
*+ bl_0_61 br_0_61 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c61
*+ bl_0_61 br_0_61 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c61
*+ bl_0_61 br_0_61 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c61
*+ bl_0_61 br_0_61 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c61
*+ bl_0_61 br_0_61 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c61
*+ bl_0_61 br_0_61 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c61
*+ bl_0_61 br_0_61 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c61
*+ bl_0_61 br_0_61 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c61
*+ bl_0_61 br_0_61 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c61
*+ bl_0_61 br_0_61 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c61
*+ bl_0_61 br_0_61 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c61
*+ bl_0_61 br_0_61 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c61
*+ bl_0_61 br_0_61 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c61
*+ bl_0_61 br_0_61 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c61
*+ bl_0_61 br_0_61 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c61
*+ bl_0_61 br_0_61 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c61
*+ bl_0_61 br_0_61 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c61
*+ bl_0_61 br_0_61 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c61
*+ bl_0_61 br_0_61 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c61
*+ bl_0_61 br_0_61 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c61
*+ bl_0_61 br_0_61 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c61
*+ bl_0_61 br_0_61 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c61
+ bl_0_61 br_0_61 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ cell_1rw
* Xbit_r1_c62
*+ bl_0_62 br_0_62 wl_0_1 vdd gnd
*+ cell_1rw
* Xbit_r2_c62
*+ bl_0_62 br_0_62 wl_0_2 vdd gnd
*+ cell_1rw
* Xbit_r3_c62
*+ bl_0_62 br_0_62 wl_0_3 vdd gnd
*+ cell_1rw
* Xbit_r4_c62
*+ bl_0_62 br_0_62 wl_0_4 vdd gnd
*+ cell_1rw
* Xbit_r5_c62
*+ bl_0_62 br_0_62 wl_0_5 vdd gnd
*+ cell_1rw
* Xbit_r6_c62
*+ bl_0_62 br_0_62 wl_0_6 vdd gnd
*+ cell_1rw
* Xbit_r7_c62
*+ bl_0_62 br_0_62 wl_0_7 vdd gnd
*+ cell_1rw
* Xbit_r8_c62
*+ bl_0_62 br_0_62 wl_0_8 vdd gnd
*+ cell_1rw
* Xbit_r9_c62
*+ bl_0_62 br_0_62 wl_0_9 vdd gnd
*+ cell_1rw
* Xbit_r10_c62
*+ bl_0_62 br_0_62 wl_0_10 vdd gnd
*+ cell_1rw
* Xbit_r11_c62
*+ bl_0_62 br_0_62 wl_0_11 vdd gnd
*+ cell_1rw
* Xbit_r12_c62
*+ bl_0_62 br_0_62 wl_0_12 vdd gnd
*+ cell_1rw
* Xbit_r13_c62
*+ bl_0_62 br_0_62 wl_0_13 vdd gnd
*+ cell_1rw
* Xbit_r14_c62
*+ bl_0_62 br_0_62 wl_0_14 vdd gnd
*+ cell_1rw
* Xbit_r15_c62
*+ bl_0_62 br_0_62 wl_0_15 vdd gnd
*+ cell_1rw
* Xbit_r16_c62
*+ bl_0_62 br_0_62 wl_0_16 vdd gnd
*+ cell_1rw
* Xbit_r17_c62
*+ bl_0_62 br_0_62 wl_0_17 vdd gnd
*+ cell_1rw
* Xbit_r18_c62
*+ bl_0_62 br_0_62 wl_0_18 vdd gnd
*+ cell_1rw
* Xbit_r19_c62
*+ bl_0_62 br_0_62 wl_0_19 vdd gnd
*+ cell_1rw
* Xbit_r20_c62
*+ bl_0_62 br_0_62 wl_0_20 vdd gnd
*+ cell_1rw
* Xbit_r21_c62
*+ bl_0_62 br_0_62 wl_0_21 vdd gnd
*+ cell_1rw
* Xbit_r22_c62
*+ bl_0_62 br_0_62 wl_0_22 vdd gnd
*+ cell_1rw
* Xbit_r23_c62
*+ bl_0_62 br_0_62 wl_0_23 vdd gnd
*+ cell_1rw
* Xbit_r24_c62
*+ bl_0_62 br_0_62 wl_0_24 vdd gnd
*+ cell_1rw
* Xbit_r25_c62
*+ bl_0_62 br_0_62 wl_0_25 vdd gnd
*+ cell_1rw
* Xbit_r26_c62
*+ bl_0_62 br_0_62 wl_0_26 vdd gnd
*+ cell_1rw
* Xbit_r27_c62
*+ bl_0_62 br_0_62 wl_0_27 vdd gnd
*+ cell_1rw
* Xbit_r28_c62
*+ bl_0_62 br_0_62 wl_0_28 vdd gnd
*+ cell_1rw
* Xbit_r29_c62
*+ bl_0_62 br_0_62 wl_0_29 vdd gnd
*+ cell_1rw
* Xbit_r30_c62
*+ bl_0_62 br_0_62 wl_0_30 vdd gnd
*+ cell_1rw
Xbit_r31_c62
+ bl_0_62 br_0_62 wl_0_31 vdd gnd
+ cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ cell_1rw
Xbit_r1_c63
+ bl_0_63 br_0_63 wl_0_1 vdd gnd
+ cell_1rw
Xbit_r2_c63
+ bl_0_63 br_0_63 wl_0_2 vdd gnd
+ cell_1rw
Xbit_r3_c63
+ bl_0_63 br_0_63 wl_0_3 vdd gnd
+ cell_1rw
Xbit_r4_c63
+ bl_0_63 br_0_63 wl_0_4 vdd gnd
+ cell_1rw
Xbit_r5_c63
+ bl_0_63 br_0_63 wl_0_5 vdd gnd
+ cell_1rw
Xbit_r6_c63
+ bl_0_63 br_0_63 wl_0_6 vdd gnd
+ cell_1rw
Xbit_r7_c63
+ bl_0_63 br_0_63 wl_0_7 vdd gnd
+ cell_1rw
Xbit_r8_c63
+ bl_0_63 br_0_63 wl_0_8 vdd gnd
+ cell_1rw
Xbit_r9_c63
+ bl_0_63 br_0_63 wl_0_9 vdd gnd
+ cell_1rw
Xbit_r10_c63
+ bl_0_63 br_0_63 wl_0_10 vdd gnd
+ cell_1rw
Xbit_r11_c63
+ bl_0_63 br_0_63 wl_0_11 vdd gnd
+ cell_1rw
Xbit_r12_c63
+ bl_0_63 br_0_63 wl_0_12 vdd gnd
+ cell_1rw
Xbit_r13_c63
+ bl_0_63 br_0_63 wl_0_13 vdd gnd
+ cell_1rw
Xbit_r14_c63
+ bl_0_63 br_0_63 wl_0_14 vdd gnd
+ cell_1rw
Xbit_r15_c63
+ bl_0_63 br_0_63 wl_0_15 vdd gnd
+ cell_1rw
Xbit_r16_c63
+ bl_0_63 br_0_63 wl_0_16 vdd gnd
+ cell_1rw
Xbit_r17_c63
+ bl_0_63 br_0_63 wl_0_17 vdd gnd
+ cell_1rw
Xbit_r18_c63
+ bl_0_63 br_0_63 wl_0_18 vdd gnd
+ cell_1rw
Xbit_r19_c63
+ bl_0_63 br_0_63 wl_0_19 vdd gnd
+ cell_1rw
Xbit_r20_c63
+ bl_0_63 br_0_63 wl_0_20 vdd gnd
+ cell_1rw
Xbit_r21_c63
+ bl_0_63 br_0_63 wl_0_21 vdd gnd
+ cell_1rw
Xbit_r22_c63
+ bl_0_63 br_0_63 wl_0_22 vdd gnd
+ cell_1rw
Xbit_r23_c63
+ bl_0_63 br_0_63 wl_0_23 vdd gnd
+ cell_1rw
Xbit_r24_c63
+ bl_0_63 br_0_63 wl_0_24 vdd gnd
+ cell_1rw
Xbit_r25_c63
+ bl_0_63 br_0_63 wl_0_25 vdd gnd
+ cell_1rw
Xbit_r26_c63
+ bl_0_63 br_0_63 wl_0_26 vdd gnd
+ cell_1rw
Xbit_r27_c63
+ bl_0_63 br_0_63 wl_0_27 vdd gnd
+ cell_1rw
Xbit_r28_c63
+ bl_0_63 br_0_63 wl_0_28 vdd gnd
+ cell_1rw
Xbit_r29_c63
+ bl_0_63 br_0_63 wl_0_29 vdd gnd
+ cell_1rw
Xbit_r30_c63
+ bl_0_63 br_0_63 wl_0_30 vdd gnd
+ cell_1rw
Xbit_r31_c63
+ bl_0_63 br_0_63 wl_0_31 vdd gnd
+ cell_1rw
.ENDS scn4m_subm_256x8_bitcell_array

.SUBCKT scn4m_subm_256x8_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 rbl_wl_0_0 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 vdd gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* POWER : vdd 
* GROUND: gnd 
* rows: 32 cols: 64
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xbitcell_array
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 vdd gnd
+ scn4m_subm_256x8_bitcell_array
Xreplica_col_0
+ rbl_bl_0_0 rbl_br_0_0 rbl_wl_0_0 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4
+ wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13
+ wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21
+ wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29
+ wl_0_30 wl_0_31 vdd gnd
+ scn4m_subm_256x8_replica_column
Xdummy_row_0
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 rbl_wl_0_0 vdd gnd
+ scn4m_subm_256x8_dummy_array
.ENDS scn4m_subm_256x8_replica_bitcell_array

.SUBCKT scn4m_subm_256x8_dummy_array_1
+ bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3 br_0_3 bl_0_4 br_0_4
+ bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8 br_0_8 bl_0_9 br_0_9
+ bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12 bl_0_13 br_0_13
+ bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16 bl_0_17 br_0_17
+ bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20 bl_0_21 br_0_21
+ bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24 bl_0_25 br_0_25
+ bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28 bl_0_29 br_0_29
+ bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32 bl_0_33 br_0_33
+ bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36 bl_0_37 br_0_37
+ bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40 bl_0_41 br_0_41
+ bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44 bl_0_45 br_0_45
+ bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48 bl_0_49 br_0_49
+ bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52 bl_0_53 br_0_53
+ bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56 bl_0_57 br_0_57
+ bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60 bl_0_61 br_0_61
+ bl_0_62 br_0_62 bl_0_63 br_0_63 bl_0_64 br_0_64 wl_0_0 vdd gnd
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INOUT : bl_0_64 
* INOUT : br_0_64 
* INPUT : wl_0_0 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_0_0 br_0_0 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c1
+ bl_0_1 br_0_1 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c2
+ bl_0_2 br_0_2 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c3
+ bl_0_3 br_0_3 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c4
+ bl_0_4 br_0_4 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c5
+ bl_0_5 br_0_5 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c6
+ bl_0_6 br_0_6 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c7
+ bl_0_7 br_0_7 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c8
+ bl_0_8 br_0_8 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c9
+ bl_0_9 br_0_9 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c10
+ bl_0_10 br_0_10 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c11
+ bl_0_11 br_0_11 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c12
+ bl_0_12 br_0_12 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c13
+ bl_0_13 br_0_13 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c14
+ bl_0_14 br_0_14 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c15
+ bl_0_15 br_0_15 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c16
+ bl_0_16 br_0_16 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c17
+ bl_0_17 br_0_17 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c18
+ bl_0_18 br_0_18 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c19
+ bl_0_19 br_0_19 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c20
+ bl_0_20 br_0_20 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c21
+ bl_0_21 br_0_21 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c22
+ bl_0_22 br_0_22 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c23
+ bl_0_23 br_0_23 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c24
+ bl_0_24 br_0_24 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c25
+ bl_0_25 br_0_25 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c26
+ bl_0_26 br_0_26 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c27
+ bl_0_27 br_0_27 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c28
+ bl_0_28 br_0_28 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c29
+ bl_0_29 br_0_29 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c30
+ bl_0_30 br_0_30 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c31
+ bl_0_31 br_0_31 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c32
+ bl_0_32 br_0_32 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c33
+ bl_0_33 br_0_33 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c34
+ bl_0_34 br_0_34 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c35
+ bl_0_35 br_0_35 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c36
+ bl_0_36 br_0_36 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c37
+ bl_0_37 br_0_37 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c38
+ bl_0_38 br_0_38 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c39
+ bl_0_39 br_0_39 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c40
+ bl_0_40 br_0_40 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c41
+ bl_0_41 br_0_41 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c42
+ bl_0_42 br_0_42 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c43
+ bl_0_43 br_0_43 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c44
+ bl_0_44 br_0_44 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c45
+ bl_0_45 br_0_45 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c46
+ bl_0_46 br_0_46 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c47
+ bl_0_47 br_0_47 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c48
+ bl_0_48 br_0_48 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c49
+ bl_0_49 br_0_49 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c50
+ bl_0_50 br_0_50 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c51
+ bl_0_51 br_0_51 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c52
+ bl_0_52 br_0_52 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c53
+ bl_0_53 br_0_53 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c54
+ bl_0_54 br_0_54 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c55
+ bl_0_55 br_0_55 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c56
+ bl_0_56 br_0_56 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c57
+ bl_0_57 br_0_57 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c58
+ bl_0_58 br_0_58 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c59
+ bl_0_59 br_0_59 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c60
+ bl_0_60 br_0_60 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c61
+ bl_0_61 br_0_61 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c62
+ bl_0_62 br_0_62 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c63
+ bl_0_63 br_0_63 wl_0_0 vdd gnd
+ dummy_cell_1rw
Xbit_r0_c64
+ bl_0_64 br_0_64 wl_0_0 vdd gnd
+ dummy_cell_1rw
.ENDS scn4m_subm_256x8_dummy_array_1

.SUBCKT scn4m_subm_256x8_capped_replica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 rbl_wl_0_0 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 vdd gnd
* INOUT : rbl_bl_0_0 
* INOUT : rbl_br_0_0 
* INOUT : bl_0_0 
* INOUT : br_0_0 
* INOUT : bl_0_1 
* INOUT : br_0_1 
* INOUT : bl_0_2 
* INOUT : br_0_2 
* INOUT : bl_0_3 
* INOUT : br_0_3 
* INOUT : bl_0_4 
* INOUT : br_0_4 
* INOUT : bl_0_5 
* INOUT : br_0_5 
* INOUT : bl_0_6 
* INOUT : br_0_6 
* INOUT : bl_0_7 
* INOUT : br_0_7 
* INOUT : bl_0_8 
* INOUT : br_0_8 
* INOUT : bl_0_9 
* INOUT : br_0_9 
* INOUT : bl_0_10 
* INOUT : br_0_10 
* INOUT : bl_0_11 
* INOUT : br_0_11 
* INOUT : bl_0_12 
* INOUT : br_0_12 
* INOUT : bl_0_13 
* INOUT : br_0_13 
* INOUT : bl_0_14 
* INOUT : br_0_14 
* INOUT : bl_0_15 
* INOUT : br_0_15 
* INOUT : bl_0_16 
* INOUT : br_0_16 
* INOUT : bl_0_17 
* INOUT : br_0_17 
* INOUT : bl_0_18 
* INOUT : br_0_18 
* INOUT : bl_0_19 
* INOUT : br_0_19 
* INOUT : bl_0_20 
* INOUT : br_0_20 
* INOUT : bl_0_21 
* INOUT : br_0_21 
* INOUT : bl_0_22 
* INOUT : br_0_22 
* INOUT : bl_0_23 
* INOUT : br_0_23 
* INOUT : bl_0_24 
* INOUT : br_0_24 
* INOUT : bl_0_25 
* INOUT : br_0_25 
* INOUT : bl_0_26 
* INOUT : br_0_26 
* INOUT : bl_0_27 
* INOUT : br_0_27 
* INOUT : bl_0_28 
* INOUT : br_0_28 
* INOUT : bl_0_29 
* INOUT : br_0_29 
* INOUT : bl_0_30 
* INOUT : br_0_30 
* INOUT : bl_0_31 
* INOUT : br_0_31 
* INOUT : bl_0_32 
* INOUT : br_0_32 
* INOUT : bl_0_33 
* INOUT : br_0_33 
* INOUT : bl_0_34 
* INOUT : br_0_34 
* INOUT : bl_0_35 
* INOUT : br_0_35 
* INOUT : bl_0_36 
* INOUT : br_0_36 
* INOUT : bl_0_37 
* INOUT : br_0_37 
* INOUT : bl_0_38 
* INOUT : br_0_38 
* INOUT : bl_0_39 
* INOUT : br_0_39 
* INOUT : bl_0_40 
* INOUT : br_0_40 
* INOUT : bl_0_41 
* INOUT : br_0_41 
* INOUT : bl_0_42 
* INOUT : br_0_42 
* INOUT : bl_0_43 
* INOUT : br_0_43 
* INOUT : bl_0_44 
* INOUT : br_0_44 
* INOUT : bl_0_45 
* INOUT : br_0_45 
* INOUT : bl_0_46 
* INOUT : br_0_46 
* INOUT : bl_0_47 
* INOUT : br_0_47 
* INOUT : bl_0_48 
* INOUT : br_0_48 
* INOUT : bl_0_49 
* INOUT : br_0_49 
* INOUT : bl_0_50 
* INOUT : br_0_50 
* INOUT : bl_0_51 
* INOUT : br_0_51 
* INOUT : bl_0_52 
* INOUT : br_0_52 
* INOUT : bl_0_53 
* INOUT : br_0_53 
* INOUT : bl_0_54 
* INOUT : br_0_54 
* INOUT : bl_0_55 
* INOUT : br_0_55 
* INOUT : bl_0_56 
* INOUT : br_0_56 
* INOUT : bl_0_57 
* INOUT : br_0_57 
* INOUT : bl_0_58 
* INOUT : br_0_58 
* INOUT : bl_0_59 
* INOUT : br_0_59 
* INOUT : bl_0_60 
* INOUT : br_0_60 
* INOUT : bl_0_61 
* INOUT : br_0_61 
* INOUT : bl_0_62 
* INOUT : br_0_62 
* INOUT : bl_0_63 
* INOUT : br_0_63 
* INPUT : rbl_wl_0_0 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* POWER : vdd 
* GROUND: gnd 
* rows: 32 cols: 64
* rbl: [1, 0] left_rbl: [0] right_rbl: []
Xreplica_bitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 rbl_wl_0_0 wl_0_0
+ wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 vdd gnd
+ scn4m_subm_256x8_replica_bitcell_array
Xdummy_row_bot
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 gnd vdd gnd
+ scn4m_subm_256x8_dummy_array_1
Xdummy_row_top
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 gnd vdd gnd
+ scn4m_subm_256x8_dummy_array_0
Xdummy_col_left
+ dummy_left_bl_0_0 dummy_left_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 gnd vdd gnd
+ scn4m_subm_256x8_dummy_array_2
Xdummy_col_right
+ dummy_right_bl_0_0 dummy_right_br_0_0 gnd rbl_wl_0_0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 gnd vdd gnd
+ scn4m_subm_256x8_dummy_array_3
.ENDS scn4m_subm_256x8_capped_replica_bitcell_array

.SUBCKT scn4m_subm_256x8_pdriver
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1]
Xbuf_inv1
+ A Z vdd gnd
+ scn4m_subm_256x8_pinv_1
.ENDS scn4m_subm_256x8_pdriver

.SUBCKT scn4m_subm_256x8_pand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_nand
+ A B C zb_int vdd gnd
+ scn4m_subm_256x8_pnand3_0
Xpand3_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pdriver
.ENDS scn4m_subm_256x8_pand3

.SUBCKT scn4m_subm_256x8_hierarchical_predecode3x8_0
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ scn4m_subm_256x8_pinv_2
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ scn4m_subm_256x8_pinv_2
Xpre_inv_2
+ in_2 inbar_2 vdd gnd
+ scn4m_subm_256x8_pinv_2
XXpre3x8_and_0
+ inbar_0 inbar_1 inbar_2 out_0 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_1
+ in_0 inbar_1 inbar_2 out_1 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_2
+ inbar_0 in_1 inbar_2 out_2 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_3
+ in_0 in_1 inbar_2 out_3 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_4
+ inbar_0 inbar_1 in_2 out_4 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_5
+ in_0 inbar_1 in_2 out_5 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_6
+ inbar_0 in_1 in_2 out_6 vdd gnd
+ scn4m_subm_256x8_pand3
XXpre3x8_and_7
+ in_0 in_1 in_2 out_7 vdd gnd
+ scn4m_subm_256x8_pand3
.ENDS scn4m_subm_256x8_hierarchical_predecode3x8_0

.SUBCKT scn4m_subm_256x8_column_decoder
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xcolumn_decoder
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
+ scn4m_subm_256x8_hierarchical_predecode3x8_0
.ENDS scn4m_subm_256x8_column_decoder

* spice ptx M{0} {1} p m=8 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p

* spice ptx M{0} {1} n m=8 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p

.SUBCKT scn4m_subm_256x8_pinv_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 16
Mpinv_pmos Z A vdd vdd p m=8 w=3.2u l=0.4u pd=7.20u ps=7.20u as=3.20p ad=3.20p
Mpinv_nmos Z A gnd gnd n m=8 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pinv_0

.SUBCKT scn4m_subm_256x8_pnand2
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand2_pmos1 vdd A Z vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pnand2

.SUBCKT scn4m_subm_256x8_and2_dec_0
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 16
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ scn4m_subm_256x8_pnand2
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pinv_0
.ENDS scn4m_subm_256x8_and2_dec_0

.SUBCKT scn4m_subm_256x8_pinv
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpinv_pmos Z A vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpinv_nmos Z A gnd gnd n m=1 w=0.8u l=0.4u pd=2.40u ps=2.40u as=0.80p ad=0.80p
.ENDS scn4m_subm_256x8_pinv

.SUBCKT scn4m_subm_256x8_and2_dec
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand2_dec_nand
+ A B zb_int vdd gnd
+ scn4m_subm_256x8_pnand2
Xpand2_dec_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pinv
.ENDS scn4m_subm_256x8_and2_dec

.SUBCKT scn4m_subm_256x8_pnand3
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Mpnand3_pmos1 vdd A Z vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=1.6u l=0.4u pd=4.00u ps=4.00u as=1.60p ad=1.60p
.ENDS scn4m_subm_256x8_pnand3

.SUBCKT scn4m_subm_256x8_and3_dec
+ A B C Z vdd gnd
* INPUT : A 
* INPUT : B 
* INPUT : C 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* size: 1
Xpand3_dec_nand
+ A B C zb_int vdd gnd
+ scn4m_subm_256x8_pnand3
Xpand3_dec_inv
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pinv
.ENDS scn4m_subm_256x8_and3_dec

.SUBCKT scn4m_subm_256x8_hierarchical_predecode3x8
+ in_0 in_1 in_2 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ scn4m_subm_256x8_pinv
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ scn4m_subm_256x8_pinv
Xpre_inv_2
+ in_2 inbar_2 vdd gnd
+ scn4m_subm_256x8_pinv
XXpre3x8_and_0
+ inbar_0 inbar_1 inbar_2 out_0 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_1
+ in_0 inbar_1 inbar_2 out_1 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_2
+ inbar_0 in_1 inbar_2 out_2 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_3
+ in_0 in_1 inbar_2 out_3 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_4
+ inbar_0 inbar_1 in_2 out_4 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_5
+ in_0 inbar_1 in_2 out_5 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_6
+ inbar_0 in_1 in_2 out_6 vdd gnd
+ scn4m_subm_256x8_and3_dec
XXpre3x8_and_7
+ in_0 in_1 in_2 out_7 vdd gnd
+ scn4m_subm_256x8_and3_dec
.ENDS scn4m_subm_256x8_hierarchical_predecode3x8

.SUBCKT scn4m_subm_256x8_hierarchical_predecode2x4
+ in_0 in_1 out_0 out_1 out_2 out_3 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* POWER : vdd 
* GROUND: gnd 
Xpre_inv_0
+ in_0 inbar_0 vdd gnd
+ scn4m_subm_256x8_pinv
Xpre_inv_1
+ in_1 inbar_1 vdd gnd
+ scn4m_subm_256x8_pinv
XXpre2x4_and_0
+ inbar_0 inbar_1 out_0 vdd gnd
+ scn4m_subm_256x8_and2_dec
XXpre2x4_and_1
+ in_0 inbar_1 out_1 vdd gnd
+ scn4m_subm_256x8_and2_dec
XXpre2x4_and_2
+ inbar_0 in_1 out_2 vdd gnd
+ scn4m_subm_256x8_and2_dec
XXpre2x4_and_3
+ in_0 in_1 out_3 vdd gnd
+ scn4m_subm_256x8_and2_dec
.ENDS scn4m_subm_256x8_hierarchical_predecode2x4

.SUBCKT scn4m_subm_256x8_hierarchical_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 decode_0 decode_1 decode_2 decode_3
+ decode_4 decode_5 decode_6 decode_7 decode_8 decode_9 decode_10
+ decode_11 decode_12 decode_13 decode_14 decode_15 decode_16 decode_17
+ decode_18 decode_19 decode_20 decode_21 decode_22 decode_23 decode_24
+ decode_25 decode_26 decode_27 decode_28 decode_29 decode_30 decode_31
+ vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* OUTPUT: decode_0 
* OUTPUT: decode_1 
* OUTPUT: decode_2 
* OUTPUT: decode_3 
* OUTPUT: decode_4 
* OUTPUT: decode_5 
* OUTPUT: decode_6 
* OUTPUT: decode_7 
* OUTPUT: decode_8 
* OUTPUT: decode_9 
* OUTPUT: decode_10 
* OUTPUT: decode_11 
* OUTPUT: decode_12 
* OUTPUT: decode_13 
* OUTPUT: decode_14 
* OUTPUT: decode_15 
* OUTPUT: decode_16 
* OUTPUT: decode_17 
* OUTPUT: decode_18 
* OUTPUT: decode_19 
* OUTPUT: decode_20 
* OUTPUT: decode_21 
* OUTPUT: decode_22 
* OUTPUT: decode_23 
* OUTPUT: decode_24 
* OUTPUT: decode_25 
* OUTPUT: decode_26 
* OUTPUT: decode_27 
* OUTPUT: decode_28 
* OUTPUT: decode_29 
* OUTPUT: decode_30 
* OUTPUT: decode_31 
* POWER : vdd 
* GROUND: gnd 
Xpre_0
+ addr_0 addr_1 out_0 out_1 out_2 out_3 vdd gnd
+ scn4m_subm_256x8_hierarchical_predecode2x4
Xpre3x8_0
+ addr_2 addr_3 addr_4 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11
+ vdd gnd
+ scn4m_subm_256x8_hierarchical_predecode3x8
XDEC_AND_0
+ out_0 out_4 decode_0 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_4
+ out_0 out_5 decode_4 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_8
+ out_0 out_6 decode_8 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_12
+ out_0 out_7 decode_12 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_16
+ out_0 out_8 decode_16 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_20
+ out_0 out_9 decode_20 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_24
+ out_0 out_10 decode_24 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_28
+ out_0 out_11 decode_28 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_1
+ out_1 out_4 decode_1 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_5
+ out_1 out_5 decode_5 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_9
+ out_1 out_6 decode_9 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_13
+ out_1 out_7 decode_13 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_17
+ out_1 out_8 decode_17 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_21
+ out_1 out_9 decode_21 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_25
+ out_1 out_10 decode_25 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_29
+ out_1 out_11 decode_29 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_2
+ out_2 out_4 decode_2 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_6
+ out_2 out_5 decode_6 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_10
+ out_2 out_6 decode_10 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_14
+ out_2 out_7 decode_14 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_18
+ out_2 out_8 decode_18 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_22
+ out_2 out_9 decode_22 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_26
+ out_2 out_10 decode_26 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_30
+ out_2 out_11 decode_30 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_3
+ out_3 out_4 decode_3 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_7
+ out_3 out_5 decode_7 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_11
+ out_3 out_6 decode_11 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_15
+ out_3 out_7 decode_15 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_19
+ out_3 out_8 decode_19 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_23
+ out_3 out_9 decode_23 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_27
+ out_3 out_10 decode_27 vdd gnd
+ scn4m_subm_256x8_and2_dec
XDEC_AND_31
+ out_3 out_11 decode_31 vdd gnd
+ scn4m_subm_256x8_and2_dec
.ENDS scn4m_subm_256x8_hierarchical_decoder

.SUBCKT scn4m_subm_256x8_wordline_driver
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* cols: 64
Xwld_nand
+ A B zb_int vdd gnd
+ scn4m_subm_256x8_pnand2
Xwl_driver
+ zb_int Z vdd gnd
+ scn4m_subm_256x8_pinv_0
.ENDS scn4m_subm_256x8_wordline_driver

.SUBCKT scn4m_subm_256x8_wordline_driver_array
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23
+ in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 wl_0 wl_1 wl_2 wl_3
+ wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 en vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* INPUT : en 
* POWER : vdd 
* GROUND: gnd 
* rows: 32 cols: 64
Xwl_driver_and0
+ in_0 en wl_0 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and1
+ in_1 en wl_1 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and2
+ in_2 en wl_2 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and3
+ in_3 en wl_3 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and4
+ in_4 en wl_4 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and5
+ in_5 en wl_5 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and6
+ in_6 en wl_6 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and7
+ in_7 en wl_7 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and8
+ in_8 en wl_8 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and9
+ in_9 en wl_9 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and10
+ in_10 en wl_10 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and11
+ in_11 en wl_11 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and12
+ in_12 en wl_12 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and13
+ in_13 en wl_13 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and14
+ in_14 en wl_14 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and15
+ in_15 en wl_15 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and16
+ in_16 en wl_16 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and17
+ in_17 en wl_17 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and18
+ in_18 en wl_18 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and19
+ in_19 en wl_19 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and20
+ in_20 en wl_20 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and21
+ in_21 en wl_21 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and22
+ in_22 en wl_22 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and23
+ in_23 en wl_23 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and24
+ in_24 en wl_24 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and25
+ in_25 en wl_25 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and26
+ in_26 en wl_26 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and27
+ in_27 en wl_27 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and28
+ in_28 en wl_28 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and29
+ in_29 en wl_29 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and30
+ in_30 en wl_30 vdd gnd
+ scn4m_subm_256x8_wordline_driver
Xwl_driver_and31
+ in_31 en wl_31 vdd gnd
+ scn4m_subm_256x8_wordline_driver
.ENDS scn4m_subm_256x8_wordline_driver_array

.SUBCKT scn4m_subm_256x8_port_address
+ addr_0 addr_1 addr_2 addr_3 addr_4 wl_en wl_0 wl_1 wl_2 wl_3 wl_4 wl_5
+ wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17
+ wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28
+ wl_29 wl_30 wl_31 rbl_wl vdd gnd
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : wl_en 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: rbl_wl 
* POWER : vdd 
* GROUND: gnd 
Xrow_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 dec_out_0 dec_out_1 dec_out_2
+ dec_out_3 dec_out_4 dec_out_5 dec_out_6 dec_out_7 dec_out_8 dec_out_9
+ dec_out_10 dec_out_11 dec_out_12 dec_out_13 dec_out_14 dec_out_15
+ dec_out_16 dec_out_17 dec_out_18 dec_out_19 dec_out_20 dec_out_21
+ dec_out_22 dec_out_23 dec_out_24 dec_out_25 dec_out_26 dec_out_27
+ dec_out_28 dec_out_29 dec_out_30 dec_out_31 vdd gnd
+ scn4m_subm_256x8_hierarchical_decoder
Xwordline_driver
+ dec_out_0 dec_out_1 dec_out_2 dec_out_3 dec_out_4 dec_out_5 dec_out_6
+ dec_out_7 dec_out_8 dec_out_9 dec_out_10 dec_out_11 dec_out_12
+ dec_out_13 dec_out_14 dec_out_15 dec_out_16 dec_out_17 dec_out_18
+ dec_out_19 dec_out_20 dec_out_21 dec_out_22 dec_out_23 dec_out_24
+ dec_out_25 dec_out_26 dec_out_27 dec_out_28 dec_out_29 dec_out_30
+ dec_out_31 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10
+ wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21
+ wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31 wl_en vdd
+ gnd
+ scn4m_subm_256x8_wordline_driver_array
Xrbl_driver
+ wl_en vdd rbl_wl vdd gnd
+ scn4m_subm_256x8_and2_dec_0
.ENDS scn4m_subm_256x8_port_address

.SUBCKT scn4m_subm_256x8_bank
+ dout0_0 dout0_1 dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7
+ rbl_bl_0_0 din0_0 din0_1 din0_2 din0_3 din0_4 din0_5 din0_6 din0_7
+ addr0_0 addr0_1 addr0_2 addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 s_en0
+ p_en_bar0 w_en0 wl_en0 vdd gnd
* OUTPUT: dout0_0 
* OUTPUT: dout0_1 
* OUTPUT: dout0_2 
* OUTPUT: dout0_3 
* OUTPUT: dout0_4 
* OUTPUT: dout0_5 
* OUTPUT: dout0_6 
* OUTPUT: dout0_7 
* OUTPUT: rbl_bl_0_0 
* INPUT : din0_0 
* INPUT : din0_1 
* INPUT : din0_2 
* INPUT : din0_3 
* INPUT : din0_4 
* INPUT : din0_5 
* INPUT : din0_6 
* INPUT : din0_7 
* INPUT : addr0_0 
* INPUT : addr0_1 
* INPUT : addr0_2 
* INPUT : addr0_3 
* INPUT : addr0_4 
* INPUT : addr0_5 
* INPUT : addr0_6 
* INPUT : addr0_7 
* INPUT : s_en0 
* INPUT : p_en_bar0 
* INPUT : w_en0 
* INPUT : wl_en0 
* POWER : vdd 
* GROUND: gnd 
Xbitcell_array
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 rbl_wl0 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18
+ wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26
+ wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 vdd gnd
+ scn4m_subm_256x8_capped_replica_bitcell_array
Xport_data0
+ rbl_bl_0_0 rbl_br_0_0 bl_0_0 br_0_0 bl_0_1 br_0_1 bl_0_2 br_0_2 bl_0_3
+ br_0_3 bl_0_4 br_0_4 bl_0_5 br_0_5 bl_0_6 br_0_6 bl_0_7 br_0_7 bl_0_8
+ br_0_8 bl_0_9 br_0_9 bl_0_10 br_0_10 bl_0_11 br_0_11 bl_0_12 br_0_12
+ bl_0_13 br_0_13 bl_0_14 br_0_14 bl_0_15 br_0_15 bl_0_16 br_0_16
+ bl_0_17 br_0_17 bl_0_18 br_0_18 bl_0_19 br_0_19 bl_0_20 br_0_20
+ bl_0_21 br_0_21 bl_0_22 br_0_22 bl_0_23 br_0_23 bl_0_24 br_0_24
+ bl_0_25 br_0_25 bl_0_26 br_0_26 bl_0_27 br_0_27 bl_0_28 br_0_28
+ bl_0_29 br_0_29 bl_0_30 br_0_30 bl_0_31 br_0_31 bl_0_32 br_0_32
+ bl_0_33 br_0_33 bl_0_34 br_0_34 bl_0_35 br_0_35 bl_0_36 br_0_36
+ bl_0_37 br_0_37 bl_0_38 br_0_38 bl_0_39 br_0_39 bl_0_40 br_0_40
+ bl_0_41 br_0_41 bl_0_42 br_0_42 bl_0_43 br_0_43 bl_0_44 br_0_44
+ bl_0_45 br_0_45 bl_0_46 br_0_46 bl_0_47 br_0_47 bl_0_48 br_0_48
+ bl_0_49 br_0_49 bl_0_50 br_0_50 bl_0_51 br_0_51 bl_0_52 br_0_52
+ bl_0_53 br_0_53 bl_0_54 br_0_54 bl_0_55 br_0_55 bl_0_56 br_0_56
+ bl_0_57 br_0_57 bl_0_58 br_0_58 bl_0_59 br_0_59 bl_0_60 br_0_60
+ bl_0_61 br_0_61 bl_0_62 br_0_62 bl_0_63 br_0_63 dout0_0 dout0_1
+ dout0_2 dout0_3 dout0_4 dout0_5 dout0_6 dout0_7 din0_0 din0_1 din0_2
+ din0_3 din0_4 din0_5 din0_6 din0_7 sel0_0 sel0_1 sel0_2 sel0_3 sel0_4
+ sel0_5 sel0_6 sel0_7 s_en0 p_en_bar0 w_en0 vdd gnd
+ scn4m_subm_256x8_port_data
Xport_address0
+ addr0_3 addr0_4 addr0_5 addr0_6 addr0_7 wl_en0 wl_0_0 wl_0_1 wl_0_2
+ wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10 wl_0_11
+ wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16 wl_0_17 wl_0_18 wl_0_19
+ wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24 wl_0_25 wl_0_26 wl_0_27
+ wl_0_28 wl_0_29 wl_0_30 wl_0_31 rbl_wl0 vdd gnd
+ scn4m_subm_256x8_port_address
Xcol_address_decoder0
+ addr0_0 addr0_1 addr0_2 sel0_0 sel0_1 sel0_2 sel0_3 sel0_4 sel0_5
+ sel0_6 sel0_7 vdd gnd
+ scn4m_subm_256x8_column_decoder
.ENDS scn4m_subm_256x8_bank

.SUBCKT scn4m_subm_256x8_row_addr_dff
+ din_0 din_1 din_2 din_3 din_4 dout_0 dout_1 dout_2 dout_3 dout_4 clk
+ vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 5 cols: 1
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r1_c0
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r2_c0
+ din_2 dout_2 clk vdd gnd
+ dff
Xdff_r3_c0
+ din_3 dout_3 clk vdd gnd
+ dff
Xdff_r4_c0
+ din_4 dout_4 clk vdd gnd
+ dff
.ENDS scn4m_subm_256x8_row_addr_dff

.SUBCKT scn4m_subm_256x8_col_addr_dff
+ din_0 din_1 din_2 dout_0 dout_1 dout_2 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 3
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r0_c1
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r0_c2
+ din_2 dout_2 clk vdd gnd
+ dff
.ENDS scn4m_subm_256x8_col_addr_dff

.SUBCKT scn4m_subm_256x8_data_dff
+ din_0 din_1 din_2 din_3 din_4 din_5 din_6 din_7 dout_0 dout_1 dout_2
+ dout_3 dout_4 dout_5 dout_6 dout_7 clk vdd gnd
* INPUT : din_0 
* INPUT : din_1 
* INPUT : din_2 
* INPUT : din_3 
* INPUT : din_4 
* INPUT : din_5 
* INPUT : din_6 
* INPUT : din_7 
* OUTPUT: dout_0 
* OUTPUT: dout_1 
* OUTPUT: dout_2 
* OUTPUT: dout_3 
* OUTPUT: dout_4 
* OUTPUT: dout_5 
* OUTPUT: dout_6 
* OUTPUT: dout_7 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
* rows: 1 cols: 8
Xdff_r0_c0
+ din_0 dout_0 clk vdd gnd
+ dff
Xdff_r0_c1
+ din_1 dout_1 clk vdd gnd
+ dff
Xdff_r0_c2
+ din_2 dout_2 clk vdd gnd
+ dff
Xdff_r0_c3
+ din_3 dout_3 clk vdd gnd
+ dff
Xdff_r0_c4
+ din_4 dout_4 clk vdd gnd
+ dff
Xdff_r0_c5
+ din_5 dout_5 clk vdd gnd
+ dff
Xdff_r0_c6
+ din_6 dout_6 clk vdd gnd
+ dff
Xdff_r0_c7
+ din_7 dout_7 clk vdd gnd
+ dff
.ENDS scn4m_subm_256x8_data_dff

.SUBCKT scn4m_subm_256x8
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] csb0 web0 clk0 dout0[0] dout0[1] dout0[2] dout0[3] dout0[4]
+ dout0[5] dout0[6] dout0[7] vdd gnd
* INPUT : din0[0] 
* INPUT : din0[1] 
* INPUT : din0[2] 
* INPUT : din0[3] 
* INPUT : din0[4] 
* INPUT : din0[5] 
* INPUT : din0[6] 
* INPUT : din0[7] 
* INPUT : addr0[0] 
* INPUT : addr0[1] 
* INPUT : addr0[2] 
* INPUT : addr0[3] 
* INPUT : addr0[4] 
* INPUT : addr0[5] 
* INPUT : addr0[6] 
* INPUT : addr0[7] 
* INPUT : csb0 
* INPUT : web0 
* INPUT : clk0 
* OUTPUT: dout0[0] 
* OUTPUT: dout0[1] 
* OUTPUT: dout0[2] 
* OUTPUT: dout0[3] 
* OUTPUT: dout0[4] 
* OUTPUT: dout0[5] 
* OUTPUT: dout0[6] 
* OUTPUT: dout0[7] 
* POWER : vdd 
* GROUND: gnd 
Xbank0
+ dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5] dout0[6]
+ dout0[7] rbl_bl0 bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3
+ bank_din0_4 bank_din0_5 bank_din0_6 bank_din0_7 a0_0 a0_1 a0_2 a0_3
+ a0_4 a0_5 a0_6 a0_7 s_en0 p_en_bar0 w_en0 wl_en0 vdd gnd
+ scn4m_subm_256x8_bank
Xcontrol0
+ csb0 web0 clk0 rbl_bl0 s_en0 w_en0 p_en_bar0 wl_en0 clk_buf0 vdd gnd
+ scn4m_subm_256x8_control_logic_rw
Xrow_address0
+ addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] a0_3 a0_4 a0_5 a0_6 a0_7
+ clk_buf0 vdd gnd
+ scn4m_subm_256x8_row_addr_dff
Xcol_address0
+ addr0[0] addr0[1] addr0[2] a0_0 a0_1 a0_2 clk_buf0 vdd gnd
+ scn4m_subm_256x8_col_addr_dff
Xdata_dff0
+ din0[0] din0[1] din0[2] din0[3] din0[4] din0[5] din0[6] din0[7]
+ bank_din0_0 bank_din0_1 bank_din0_2 bank_din0_3 bank_din0_4
+ bank_din0_5 bank_din0_6 bank_din0_7 clk_buf0 vdd gnd
+ scn4m_subm_256x8_data_dff
.ENDS scn4m_subm_256x8
