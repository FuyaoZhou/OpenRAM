VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45-spice-710-128x8
   CLASS BLOCK ;
   SIZE 60.805 BY 74.485 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  26.1675 0.0 26.3075 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  29.0275 0.0 29.1675 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  31.8875 0.0 32.0275 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  34.7475 0.0 34.8875 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  37.6075 0.0 37.7475 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  40.4675 0.0 40.6075 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  43.3275 0.0 43.4675 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  46.1875 0.0 46.3275 0.14 ;
      END
   END din0[7]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  20.4475 0.0 20.5875 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  23.3075 0.0 23.4475 0.14 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 46.24 0.14 46.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 48.97 0.14 49.11 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 51.18 0.14 51.32 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 53.91 0.14 54.05 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 56.12 0.14 56.26 ;
      END
   END addr0[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 4.25 0.14 4.39 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 6.98 0.14 7.12 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.84 0.0 9.98 0.14 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.2875 0.0 33.4275 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.1075 0.0 36.2475 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  38.9275 0.0 39.0675 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  41.7475 0.0 41.8875 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.5675 0.0 44.7075 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.3875 0.0 47.5275 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.665 12.4125 60.805 12.5525 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  60.665 12.1775 60.805 12.3175 ;
      END
   END dout0[7]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 0.0 60.805 0.7 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 74.485 ;
         LAYER metal3 ;
         RECT  0.0 73.785 60.805 74.485 ;
         LAYER metal4 ;
         RECT  60.105 0.0 60.805 74.485 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 73.085 ;
         LAYER metal4 ;
         RECT  58.705 1.4 59.405 73.085 ;
         LAYER metal3 ;
         RECT  1.4 72.385 59.405 73.085 ;
         LAYER metal3 ;
         RECT  1.4 1.4 59.405 2.1 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 60.665 74.345 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 60.665 74.345 ;
   LAYER  metal3 ;
      RECT  0.28 46.1 60.665 46.52 ;
      RECT  0.14 46.52 0.28 48.83 ;
      RECT  0.14 49.25 0.28 51.04 ;
      RECT  0.14 51.46 0.28 53.77 ;
      RECT  0.14 54.19 0.28 55.98 ;
      RECT  0.14 4.53 0.28 6.84 ;
      RECT  0.14 7.26 0.28 46.1 ;
      RECT  0.28 12.2725 60.525 12.6925 ;
      RECT  0.28 12.6925 60.525 46.1 ;
      RECT  60.525 12.6925 60.665 46.1 ;
      RECT  0.14 0.84 0.28 4.11 ;
      RECT  60.525 0.84 60.665 12.0375 ;
      RECT  0.14 56.4 0.28 73.645 ;
      RECT  0.28 46.52 1.26 72.245 ;
      RECT  0.28 72.245 1.26 73.225 ;
      RECT  0.28 73.225 1.26 73.645 ;
      RECT  1.26 46.52 59.545 72.245 ;
      RECT  1.26 73.225 59.545 73.645 ;
      RECT  59.545 46.52 60.665 72.245 ;
      RECT  59.545 72.245 60.665 73.225 ;
      RECT  59.545 73.225 60.665 73.645 ;
      RECT  0.28 0.84 1.26 1.26 ;
      RECT  0.28 1.26 1.26 2.24 ;
      RECT  0.28 2.24 1.26 12.2725 ;
      RECT  1.26 0.84 59.545 1.26 ;
      RECT  1.26 2.24 59.545 12.2725 ;
      RECT  59.545 0.84 60.525 1.26 ;
      RECT  59.545 1.26 60.525 2.24 ;
      RECT  59.545 2.24 60.525 12.2725 ;
   LAYER  metal4 ;
      RECT  25.8875 0.42 26.5875 74.345 ;
      RECT  26.5875 0.14 28.7475 0.42 ;
      RECT  29.4475 0.14 31.6075 0.42 ;
      RECT  20.8675 0.14 23.0275 0.42 ;
      RECT  23.7275 0.14 25.8875 0.42 ;
      RECT  10.26 0.14 20.1675 0.42 ;
      RECT  32.3075 0.14 33.0075 0.42 ;
      RECT  33.7075 0.14 34.4675 0.42 ;
      RECT  35.1675 0.14 35.8275 0.42 ;
      RECT  36.5275 0.14 37.3275 0.42 ;
      RECT  38.0275 0.14 38.6475 0.42 ;
      RECT  39.3475 0.14 40.1875 0.42 ;
      RECT  40.8875 0.14 41.4675 0.42 ;
      RECT  42.1675 0.14 43.0475 0.42 ;
      RECT  43.7475 0.14 44.2875 0.42 ;
      RECT  44.9875 0.14 45.9075 0.42 ;
      RECT  46.6075 0.14 47.1075 0.42 ;
      RECT  0.98 0.14 9.56 0.42 ;
      RECT  47.8075 0.14 59.825 0.42 ;
      RECT  0.98 0.42 1.12 1.12 ;
      RECT  0.98 1.12 1.12 73.365 ;
      RECT  0.98 73.365 1.12 74.345 ;
      RECT  1.12 0.42 2.38 1.12 ;
      RECT  1.12 73.365 2.38 74.345 ;
      RECT  2.38 0.42 25.8875 1.12 ;
      RECT  2.38 1.12 25.8875 73.365 ;
      RECT  2.38 73.365 25.8875 74.345 ;
      RECT  26.5875 0.42 58.425 1.12 ;
      RECT  26.5875 1.12 58.425 73.365 ;
      RECT  26.5875 73.365 58.425 74.345 ;
      RECT  58.425 0.42 59.685 1.12 ;
      RECT  58.425 73.365 59.685 74.345 ;
      RECT  59.685 0.42 59.825 1.12 ;
      RECT  59.685 1.12 59.825 73.365 ;
      RECT  59.685 73.365 59.825 74.345 ;
   END
END    freepdk45-spice-710-128x8
END    LIBRARY
